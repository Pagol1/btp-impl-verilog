`include "my_defines.vh"
`include "cla_gen_prop.v"
`include "rca.v"
`include "rcha.v"

module fxp32s_dadda(
	input clk,
	input [`FXP32S_ADDR] in_a,		// Sign-Mag
	input [`FXP32S_ADDR] in_b,		// Sign-Mag
	output [`FXP32S_ADDR] out_s,
	output out_overflow
);

	wire neg_out;
	assign neg_out = in_a[`FXP32S_SIGN] ^ in_b[`FXP32S_SIGN];
	wire [`FXP32S_ADDR] a, b;
	assign a[`FXP32S_SIGN] = 1'b0;
	assign a[`FXP32S_MAG] = in_a[`FXP32S_MAG];
	assign b[`FXP32S_SIGN] = 1'b0;
	assign b[`FXP32S_MAG] = in_b[`FXP32S_MAG];

	wire [0:0] dm_int_st0_0;
	wire [1:0] dm_int_st0_1;
	wire [2:0] dm_int_st0_2;
	wire [3:0] dm_int_st0_3;
	wire [4:0] dm_int_st0_4;
	wire [5:0] dm_int_st0_5;
	wire [6:0] dm_int_st0_6;
	wire [7:0] dm_int_st0_7;
	wire [8:0] dm_int_st0_8;
	wire [9:0] dm_int_st0_9;
	wire [10:0] dm_int_st0_10;
	wire [11:0] dm_int_st0_11;
	wire [12:0] dm_int_st0_12;
	wire [13:0] dm_int_st0_13;
	wire [14:0] dm_int_st0_14;
	wire [15:0] dm_int_st0_15;
	wire [16:0] dm_int_st0_16;
	wire [17:0] dm_int_st0_17;
	wire [18:0] dm_int_st0_18;
	wire [19:0] dm_int_st0_19;
	wire [20:0] dm_int_st0_20;
	wire [21:0] dm_int_st0_21;
	wire [22:0] dm_int_st0_22;
	wire [23:0] dm_int_st0_23;
	wire [24:0] dm_int_st0_24;
	wire [25:0] dm_int_st0_25;
	wire [26:0] dm_int_st0_26;
	wire [27:0] dm_int_st0_27;
	wire [28:0] dm_int_st0_28;
	wire [29:0] dm_int_st0_29;
	wire [30:0] dm_int_st0_30;
	wire [31:0] dm_int_st0_31;
	wire [30:0] dm_int_st0_32;
	wire [29:0] dm_int_st0_33;
	wire [28:0] dm_int_st0_34;
	wire [27:0] dm_int_st0_35;
	wire [26:0] dm_int_st0_36;
	wire [25:0] dm_int_st0_37;
	wire [24:0] dm_int_st0_38;
	wire [23:0] dm_int_st0_39;
	wire [22:0] dm_int_st0_40;
	wire [21:0] dm_int_st0_41;
	wire [20:0] dm_int_st0_42;
	wire [19:0] dm_int_st0_43;
	wire [18:0] dm_int_st0_44;
	wire [17:0] dm_int_st0_45;
	wire [16:0] dm_int_st0_46;
	wire [15:0] dm_int_st0_47;
	wire [14:0] dm_int_st0_48;
	wire [13:0] dm_int_st0_49;
	wire [12:0] dm_int_st0_50;
	wire [11:0] dm_int_st0_51;
	wire [10:0] dm_int_st0_52;
	wire [9:0] dm_int_st0_53;
	wire [8:0] dm_int_st0_54;
	wire [7:0] dm_int_st0_55;
	wire [6:0] dm_int_st0_56;
	wire [5:0] dm_int_st0_57;
	wire [4:0] dm_int_st0_58;
	wire [3:0] dm_int_st0_59;
	wire [2:0] dm_int_st0_60;
	wire [1:0] dm_int_st0_61;
	wire [0:0] dm_int_st0_62;

	assign dm_int_st0_0[0] = a[0] & b[0];
	assign dm_int_st0_1[0] = a[0] & b[1];
	assign dm_int_st0_2[0] = a[0] & b[2];
	assign dm_int_st0_3[0] = a[0] & b[3];
	assign dm_int_st0_4[0] = a[0] & b[4];
	assign dm_int_st0_5[0] = a[0] & b[5];
	assign dm_int_st0_6[0] = a[0] & b[6];
	assign dm_int_st0_7[0] = a[0] & b[7];
	assign dm_int_st0_8[0] = a[0] & b[8];
	assign dm_int_st0_9[0] = a[0] & b[9];
	assign dm_int_st0_10[0] = a[0] & b[10];
	assign dm_int_st0_11[0] = a[0] & b[11];
	assign dm_int_st0_12[0] = a[0] & b[12];
	assign dm_int_st0_13[0] = a[0] & b[13];
	assign dm_int_st0_14[0] = a[0] & b[14];
	assign dm_int_st0_15[0] = a[0] & b[15];
	assign dm_int_st0_16[0] = a[0] & b[16];
	assign dm_int_st0_17[0] = a[0] & b[17];
	assign dm_int_st0_18[0] = a[0] & b[18];
	assign dm_int_st0_19[0] = a[0] & b[19];
	assign dm_int_st0_20[0] = a[0] & b[20];
	assign dm_int_st0_21[0] = a[0] & b[21];
	assign dm_int_st0_22[0] = a[0] & b[22];
	assign dm_int_st0_23[0] = a[0] & b[23];
	assign dm_int_st0_24[0] = a[0] & b[24];
	assign dm_int_st0_25[0] = a[0] & b[25];
	assign dm_int_st0_26[0] = a[0] & b[26];
	assign dm_int_st0_27[0] = a[0] & b[27];
	assign dm_int_st0_28[0] = a[0] & b[28];
	assign dm_int_st0_29[0] = a[0] & b[29];
	assign dm_int_st0_30[0] = a[0] & b[30];
	assign dm_int_st0_31[0] = a[0] & b[31];
	assign dm_int_st0_1[1] = a[1] & b[0];
	assign dm_int_st0_2[1] = a[1] & b[1];
	assign dm_int_st0_3[1] = a[1] & b[2];
	assign dm_int_st0_4[1] = a[1] & b[3];
	assign dm_int_st0_5[1] = a[1] & b[4];
	assign dm_int_st0_6[1] = a[1] & b[5];
	assign dm_int_st0_7[1] = a[1] & b[6];
	assign dm_int_st0_8[1] = a[1] & b[7];
	assign dm_int_st0_9[1] = a[1] & b[8];
	assign dm_int_st0_10[1] = a[1] & b[9];
	assign dm_int_st0_11[1] = a[1] & b[10];
	assign dm_int_st0_12[1] = a[1] & b[11];
	assign dm_int_st0_13[1] = a[1] & b[12];
	assign dm_int_st0_14[1] = a[1] & b[13];
	assign dm_int_st0_15[1] = a[1] & b[14];
	assign dm_int_st0_16[1] = a[1] & b[15];
	assign dm_int_st0_17[1] = a[1] & b[16];
	assign dm_int_st0_18[1] = a[1] & b[17];
	assign dm_int_st0_19[1] = a[1] & b[18];
	assign dm_int_st0_20[1] = a[1] & b[19];
	assign dm_int_st0_21[1] = a[1] & b[20];
	assign dm_int_st0_22[1] = a[1] & b[21];
	assign dm_int_st0_23[1] = a[1] & b[22];
	assign dm_int_st0_24[1] = a[1] & b[23];
	assign dm_int_st0_25[1] = a[1] & b[24];
	assign dm_int_st0_26[1] = a[1] & b[25];
	assign dm_int_st0_27[1] = a[1] & b[26];
	assign dm_int_st0_28[1] = a[1] & b[27];
	assign dm_int_st0_29[1] = a[1] & b[28];
	assign dm_int_st0_30[1] = a[1] & b[29];
	assign dm_int_st0_31[1] = a[1] & b[30];
	assign dm_int_st0_32[0] = a[1] & b[31];
	assign dm_int_st0_2[2] = a[2] & b[0];
	assign dm_int_st0_3[2] = a[2] & b[1];
	assign dm_int_st0_4[2] = a[2] & b[2];
	assign dm_int_st0_5[2] = a[2] & b[3];
	assign dm_int_st0_6[2] = a[2] & b[4];
	assign dm_int_st0_7[2] = a[2] & b[5];
	assign dm_int_st0_8[2] = a[2] & b[6];
	assign dm_int_st0_9[2] = a[2] & b[7];
	assign dm_int_st0_10[2] = a[2] & b[8];
	assign dm_int_st0_11[2] = a[2] & b[9];
	assign dm_int_st0_12[2] = a[2] & b[10];
	assign dm_int_st0_13[2] = a[2] & b[11];
	assign dm_int_st0_14[2] = a[2] & b[12];
	assign dm_int_st0_15[2] = a[2] & b[13];
	assign dm_int_st0_16[2] = a[2] & b[14];
	assign dm_int_st0_17[2] = a[2] & b[15];
	assign dm_int_st0_18[2] = a[2] & b[16];
	assign dm_int_st0_19[2] = a[2] & b[17];
	assign dm_int_st0_20[2] = a[2] & b[18];
	assign dm_int_st0_21[2] = a[2] & b[19];
	assign dm_int_st0_22[2] = a[2] & b[20];
	assign dm_int_st0_23[2] = a[2] & b[21];
	assign dm_int_st0_24[2] = a[2] & b[22];
	assign dm_int_st0_25[2] = a[2] & b[23];
	assign dm_int_st0_26[2] = a[2] & b[24];
	assign dm_int_st0_27[2] = a[2] & b[25];
	assign dm_int_st0_28[2] = a[2] & b[26];
	assign dm_int_st0_29[2] = a[2] & b[27];
	assign dm_int_st0_30[2] = a[2] & b[28];
	assign dm_int_st0_31[2] = a[2] & b[29];
	assign dm_int_st0_32[1] = a[2] & b[30];
	assign dm_int_st0_33[0] = a[2] & b[31];
	assign dm_int_st0_3[3] = a[3] & b[0];
	assign dm_int_st0_4[3] = a[3] & b[1];
	assign dm_int_st0_5[3] = a[3] & b[2];
	assign dm_int_st0_6[3] = a[3] & b[3];
	assign dm_int_st0_7[3] = a[3] & b[4];
	assign dm_int_st0_8[3] = a[3] & b[5];
	assign dm_int_st0_9[3] = a[3] & b[6];
	assign dm_int_st0_10[3] = a[3] & b[7];
	assign dm_int_st0_11[3] = a[3] & b[8];
	assign dm_int_st0_12[3] = a[3] & b[9];
	assign dm_int_st0_13[3] = a[3] & b[10];
	assign dm_int_st0_14[3] = a[3] & b[11];
	assign dm_int_st0_15[3] = a[3] & b[12];
	assign dm_int_st0_16[3] = a[3] & b[13];
	assign dm_int_st0_17[3] = a[3] & b[14];
	assign dm_int_st0_18[3] = a[3] & b[15];
	assign dm_int_st0_19[3] = a[3] & b[16];
	assign dm_int_st0_20[3] = a[3] & b[17];
	assign dm_int_st0_21[3] = a[3] & b[18];
	assign dm_int_st0_22[3] = a[3] & b[19];
	assign dm_int_st0_23[3] = a[3] & b[20];
	assign dm_int_st0_24[3] = a[3] & b[21];
	assign dm_int_st0_25[3] = a[3] & b[22];
	assign dm_int_st0_26[3] = a[3] & b[23];
	assign dm_int_st0_27[3] = a[3] & b[24];
	assign dm_int_st0_28[3] = a[3] & b[25];
	assign dm_int_st0_29[3] = a[3] & b[26];
	assign dm_int_st0_30[3] = a[3] & b[27];
	assign dm_int_st0_31[3] = a[3] & b[28];
	assign dm_int_st0_32[2] = a[3] & b[29];
	assign dm_int_st0_33[1] = a[3] & b[30];
	assign dm_int_st0_34[0] = a[3] & b[31];
	assign dm_int_st0_4[4] = a[4] & b[0];
	assign dm_int_st0_5[4] = a[4] & b[1];
	assign dm_int_st0_6[4] = a[4] & b[2];
	assign dm_int_st0_7[4] = a[4] & b[3];
	assign dm_int_st0_8[4] = a[4] & b[4];
	assign dm_int_st0_9[4] = a[4] & b[5];
	assign dm_int_st0_10[4] = a[4] & b[6];
	assign dm_int_st0_11[4] = a[4] & b[7];
	assign dm_int_st0_12[4] = a[4] & b[8];
	assign dm_int_st0_13[4] = a[4] & b[9];
	assign dm_int_st0_14[4] = a[4] & b[10];
	assign dm_int_st0_15[4] = a[4] & b[11];
	assign dm_int_st0_16[4] = a[4] & b[12];
	assign dm_int_st0_17[4] = a[4] & b[13];
	assign dm_int_st0_18[4] = a[4] & b[14];
	assign dm_int_st0_19[4] = a[4] & b[15];
	assign dm_int_st0_20[4] = a[4] & b[16];
	assign dm_int_st0_21[4] = a[4] & b[17];
	assign dm_int_st0_22[4] = a[4] & b[18];
	assign dm_int_st0_23[4] = a[4] & b[19];
	assign dm_int_st0_24[4] = a[4] & b[20];
	assign dm_int_st0_25[4] = a[4] & b[21];
	assign dm_int_st0_26[4] = a[4] & b[22];
	assign dm_int_st0_27[4] = a[4] & b[23];
	assign dm_int_st0_28[4] = a[4] & b[24];
	assign dm_int_st0_29[4] = a[4] & b[25];
	assign dm_int_st0_30[4] = a[4] & b[26];
	assign dm_int_st0_31[4] = a[4] & b[27];
	assign dm_int_st0_32[3] = a[4] & b[28];
	assign dm_int_st0_33[2] = a[4] & b[29];
	assign dm_int_st0_34[1] = a[4] & b[30];
	assign dm_int_st0_35[0] = a[4] & b[31];
	assign dm_int_st0_5[5] = a[5] & b[0];
	assign dm_int_st0_6[5] = a[5] & b[1];
	assign dm_int_st0_7[5] = a[5] & b[2];
	assign dm_int_st0_8[5] = a[5] & b[3];
	assign dm_int_st0_9[5] = a[5] & b[4];
	assign dm_int_st0_10[5] = a[5] & b[5];
	assign dm_int_st0_11[5] = a[5] & b[6];
	assign dm_int_st0_12[5] = a[5] & b[7];
	assign dm_int_st0_13[5] = a[5] & b[8];
	assign dm_int_st0_14[5] = a[5] & b[9];
	assign dm_int_st0_15[5] = a[5] & b[10];
	assign dm_int_st0_16[5] = a[5] & b[11];
	assign dm_int_st0_17[5] = a[5] & b[12];
	assign dm_int_st0_18[5] = a[5] & b[13];
	assign dm_int_st0_19[5] = a[5] & b[14];
	assign dm_int_st0_20[5] = a[5] & b[15];
	assign dm_int_st0_21[5] = a[5] & b[16];
	assign dm_int_st0_22[5] = a[5] & b[17];
	assign dm_int_st0_23[5] = a[5] & b[18];
	assign dm_int_st0_24[5] = a[5] & b[19];
	assign dm_int_st0_25[5] = a[5] & b[20];
	assign dm_int_st0_26[5] = a[5] & b[21];
	assign dm_int_st0_27[5] = a[5] & b[22];
	assign dm_int_st0_28[5] = a[5] & b[23];
	assign dm_int_st0_29[5] = a[5] & b[24];
	assign dm_int_st0_30[5] = a[5] & b[25];
	assign dm_int_st0_31[5] = a[5] & b[26];
	assign dm_int_st0_32[4] = a[5] & b[27];
	assign dm_int_st0_33[3] = a[5] & b[28];
	assign dm_int_st0_34[2] = a[5] & b[29];
	assign dm_int_st0_35[1] = a[5] & b[30];
	assign dm_int_st0_36[0] = a[5] & b[31];
	assign dm_int_st0_6[6] = a[6] & b[0];
	assign dm_int_st0_7[6] = a[6] & b[1];
	assign dm_int_st0_8[6] = a[6] & b[2];
	assign dm_int_st0_9[6] = a[6] & b[3];
	assign dm_int_st0_10[6] = a[6] & b[4];
	assign dm_int_st0_11[6] = a[6] & b[5];
	assign dm_int_st0_12[6] = a[6] & b[6];
	assign dm_int_st0_13[6] = a[6] & b[7];
	assign dm_int_st0_14[6] = a[6] & b[8];
	assign dm_int_st0_15[6] = a[6] & b[9];
	assign dm_int_st0_16[6] = a[6] & b[10];
	assign dm_int_st0_17[6] = a[6] & b[11];
	assign dm_int_st0_18[6] = a[6] & b[12];
	assign dm_int_st0_19[6] = a[6] & b[13];
	assign dm_int_st0_20[6] = a[6] & b[14];
	assign dm_int_st0_21[6] = a[6] & b[15];
	assign dm_int_st0_22[6] = a[6] & b[16];
	assign dm_int_st0_23[6] = a[6] & b[17];
	assign dm_int_st0_24[6] = a[6] & b[18];
	assign dm_int_st0_25[6] = a[6] & b[19];
	assign dm_int_st0_26[6] = a[6] & b[20];
	assign dm_int_st0_27[6] = a[6] & b[21];
	assign dm_int_st0_28[6] = a[6] & b[22];
	assign dm_int_st0_29[6] = a[6] & b[23];
	assign dm_int_st0_30[6] = a[6] & b[24];
	assign dm_int_st0_31[6] = a[6] & b[25];
	assign dm_int_st0_32[5] = a[6] & b[26];
	assign dm_int_st0_33[4] = a[6] & b[27];
	assign dm_int_st0_34[3] = a[6] & b[28];
	assign dm_int_st0_35[2] = a[6] & b[29];
	assign dm_int_st0_36[1] = a[6] & b[30];
	assign dm_int_st0_37[0] = a[6] & b[31];
	assign dm_int_st0_7[7] = a[7] & b[0];
	assign dm_int_st0_8[7] = a[7] & b[1];
	assign dm_int_st0_9[7] = a[7] & b[2];
	assign dm_int_st0_10[7] = a[7] & b[3];
	assign dm_int_st0_11[7] = a[7] & b[4];
	assign dm_int_st0_12[7] = a[7] & b[5];
	assign dm_int_st0_13[7] = a[7] & b[6];
	assign dm_int_st0_14[7] = a[7] & b[7];
	assign dm_int_st0_15[7] = a[7] & b[8];
	assign dm_int_st0_16[7] = a[7] & b[9];
	assign dm_int_st0_17[7] = a[7] & b[10];
	assign dm_int_st0_18[7] = a[7] & b[11];
	assign dm_int_st0_19[7] = a[7] & b[12];
	assign dm_int_st0_20[7] = a[7] & b[13];
	assign dm_int_st0_21[7] = a[7] & b[14];
	assign dm_int_st0_22[7] = a[7] & b[15];
	assign dm_int_st0_23[7] = a[7] & b[16];
	assign dm_int_st0_24[7] = a[7] & b[17];
	assign dm_int_st0_25[7] = a[7] & b[18];
	assign dm_int_st0_26[7] = a[7] & b[19];
	assign dm_int_st0_27[7] = a[7] & b[20];
	assign dm_int_st0_28[7] = a[7] & b[21];
	assign dm_int_st0_29[7] = a[7] & b[22];
	assign dm_int_st0_30[7] = a[7] & b[23];
	assign dm_int_st0_31[7] = a[7] & b[24];
	assign dm_int_st0_32[6] = a[7] & b[25];
	assign dm_int_st0_33[5] = a[7] & b[26];
	assign dm_int_st0_34[4] = a[7] & b[27];
	assign dm_int_st0_35[3] = a[7] & b[28];
	assign dm_int_st0_36[2] = a[7] & b[29];
	assign dm_int_st0_37[1] = a[7] & b[30];
	assign dm_int_st0_38[0] = a[7] & b[31];
	assign dm_int_st0_8[8] = a[8] & b[0];
	assign dm_int_st0_9[8] = a[8] & b[1];
	assign dm_int_st0_10[8] = a[8] & b[2];
	assign dm_int_st0_11[8] = a[8] & b[3];
	assign dm_int_st0_12[8] = a[8] & b[4];
	assign dm_int_st0_13[8] = a[8] & b[5];
	assign dm_int_st0_14[8] = a[8] & b[6];
	assign dm_int_st0_15[8] = a[8] & b[7];
	assign dm_int_st0_16[8] = a[8] & b[8];
	assign dm_int_st0_17[8] = a[8] & b[9];
	assign dm_int_st0_18[8] = a[8] & b[10];
	assign dm_int_st0_19[8] = a[8] & b[11];
	assign dm_int_st0_20[8] = a[8] & b[12];
	assign dm_int_st0_21[8] = a[8] & b[13];
	assign dm_int_st0_22[8] = a[8] & b[14];
	assign dm_int_st0_23[8] = a[8] & b[15];
	assign dm_int_st0_24[8] = a[8] & b[16];
	assign dm_int_st0_25[8] = a[8] & b[17];
	assign dm_int_st0_26[8] = a[8] & b[18];
	assign dm_int_st0_27[8] = a[8] & b[19];
	assign dm_int_st0_28[8] = a[8] & b[20];
	assign dm_int_st0_29[8] = a[8] & b[21];
	assign dm_int_st0_30[8] = a[8] & b[22];
	assign dm_int_st0_31[8] = a[8] & b[23];
	assign dm_int_st0_32[7] = a[8] & b[24];
	assign dm_int_st0_33[6] = a[8] & b[25];
	assign dm_int_st0_34[5] = a[8] & b[26];
	assign dm_int_st0_35[4] = a[8] & b[27];
	assign dm_int_st0_36[3] = a[8] & b[28];
	assign dm_int_st0_37[2] = a[8] & b[29];
	assign dm_int_st0_38[1] = a[8] & b[30];
	assign dm_int_st0_39[0] = a[8] & b[31];
	assign dm_int_st0_9[9] = a[9] & b[0];
	assign dm_int_st0_10[9] = a[9] & b[1];
	assign dm_int_st0_11[9] = a[9] & b[2];
	assign dm_int_st0_12[9] = a[9] & b[3];
	assign dm_int_st0_13[9] = a[9] & b[4];
	assign dm_int_st0_14[9] = a[9] & b[5];
	assign dm_int_st0_15[9] = a[9] & b[6];
	assign dm_int_st0_16[9] = a[9] & b[7];
	assign dm_int_st0_17[9] = a[9] & b[8];
	assign dm_int_st0_18[9] = a[9] & b[9];
	assign dm_int_st0_19[9] = a[9] & b[10];
	assign dm_int_st0_20[9] = a[9] & b[11];
	assign dm_int_st0_21[9] = a[9] & b[12];
	assign dm_int_st0_22[9] = a[9] & b[13];
	assign dm_int_st0_23[9] = a[9] & b[14];
	assign dm_int_st0_24[9] = a[9] & b[15];
	assign dm_int_st0_25[9] = a[9] & b[16];
	assign dm_int_st0_26[9] = a[9] & b[17];
	assign dm_int_st0_27[9] = a[9] & b[18];
	assign dm_int_st0_28[9] = a[9] & b[19];
	assign dm_int_st0_29[9] = a[9] & b[20];
	assign dm_int_st0_30[9] = a[9] & b[21];
	assign dm_int_st0_31[9] = a[9] & b[22];
	assign dm_int_st0_32[8] = a[9] & b[23];
	assign dm_int_st0_33[7] = a[9] & b[24];
	assign dm_int_st0_34[6] = a[9] & b[25];
	assign dm_int_st0_35[5] = a[9] & b[26];
	assign dm_int_st0_36[4] = a[9] & b[27];
	assign dm_int_st0_37[3] = a[9] & b[28];
	assign dm_int_st0_38[2] = a[9] & b[29];
	assign dm_int_st0_39[1] = a[9] & b[30];
	assign dm_int_st0_40[0] = a[9] & b[31];
	assign dm_int_st0_10[10] = a[10] & b[0];
	assign dm_int_st0_11[10] = a[10] & b[1];
	assign dm_int_st0_12[10] = a[10] & b[2];
	assign dm_int_st0_13[10] = a[10] & b[3];
	assign dm_int_st0_14[10] = a[10] & b[4];
	assign dm_int_st0_15[10] = a[10] & b[5];
	assign dm_int_st0_16[10] = a[10] & b[6];
	assign dm_int_st0_17[10] = a[10] & b[7];
	assign dm_int_st0_18[10] = a[10] & b[8];
	assign dm_int_st0_19[10] = a[10] & b[9];
	assign dm_int_st0_20[10] = a[10] & b[10];
	assign dm_int_st0_21[10] = a[10] & b[11];
	assign dm_int_st0_22[10] = a[10] & b[12];
	assign dm_int_st0_23[10] = a[10] & b[13];
	assign dm_int_st0_24[10] = a[10] & b[14];
	assign dm_int_st0_25[10] = a[10] & b[15];
	assign dm_int_st0_26[10] = a[10] & b[16];
	assign dm_int_st0_27[10] = a[10] & b[17];
	assign dm_int_st0_28[10] = a[10] & b[18];
	assign dm_int_st0_29[10] = a[10] & b[19];
	assign dm_int_st0_30[10] = a[10] & b[20];
	assign dm_int_st0_31[10] = a[10] & b[21];
	assign dm_int_st0_32[9] = a[10] & b[22];
	assign dm_int_st0_33[8] = a[10] & b[23];
	assign dm_int_st0_34[7] = a[10] & b[24];
	assign dm_int_st0_35[6] = a[10] & b[25];
	assign dm_int_st0_36[5] = a[10] & b[26];
	assign dm_int_st0_37[4] = a[10] & b[27];
	assign dm_int_st0_38[3] = a[10] & b[28];
	assign dm_int_st0_39[2] = a[10] & b[29];
	assign dm_int_st0_40[1] = a[10] & b[30];
	assign dm_int_st0_41[0] = a[10] & b[31];
	assign dm_int_st0_11[11] = a[11] & b[0];
	assign dm_int_st0_12[11] = a[11] & b[1];
	assign dm_int_st0_13[11] = a[11] & b[2];
	assign dm_int_st0_14[11] = a[11] & b[3];
	assign dm_int_st0_15[11] = a[11] & b[4];
	assign dm_int_st0_16[11] = a[11] & b[5];
	assign dm_int_st0_17[11] = a[11] & b[6];
	assign dm_int_st0_18[11] = a[11] & b[7];
	assign dm_int_st0_19[11] = a[11] & b[8];
	assign dm_int_st0_20[11] = a[11] & b[9];
	assign dm_int_st0_21[11] = a[11] & b[10];
	assign dm_int_st0_22[11] = a[11] & b[11];
	assign dm_int_st0_23[11] = a[11] & b[12];
	assign dm_int_st0_24[11] = a[11] & b[13];
	assign dm_int_st0_25[11] = a[11] & b[14];
	assign dm_int_st0_26[11] = a[11] & b[15];
	assign dm_int_st0_27[11] = a[11] & b[16];
	assign dm_int_st0_28[11] = a[11] & b[17];
	assign dm_int_st0_29[11] = a[11] & b[18];
	assign dm_int_st0_30[11] = a[11] & b[19];
	assign dm_int_st0_31[11] = a[11] & b[20];
	assign dm_int_st0_32[10] = a[11] & b[21];
	assign dm_int_st0_33[9] = a[11] & b[22];
	assign dm_int_st0_34[8] = a[11] & b[23];
	assign dm_int_st0_35[7] = a[11] & b[24];
	assign dm_int_st0_36[6] = a[11] & b[25];
	assign dm_int_st0_37[5] = a[11] & b[26];
	assign dm_int_st0_38[4] = a[11] & b[27];
	assign dm_int_st0_39[3] = a[11] & b[28];
	assign dm_int_st0_40[2] = a[11] & b[29];
	assign dm_int_st0_41[1] = a[11] & b[30];
	assign dm_int_st0_42[0] = a[11] & b[31];
	assign dm_int_st0_12[12] = a[12] & b[0];
	assign dm_int_st0_13[12] = a[12] & b[1];
	assign dm_int_st0_14[12] = a[12] & b[2];
	assign dm_int_st0_15[12] = a[12] & b[3];
	assign dm_int_st0_16[12] = a[12] & b[4];
	assign dm_int_st0_17[12] = a[12] & b[5];
	assign dm_int_st0_18[12] = a[12] & b[6];
	assign dm_int_st0_19[12] = a[12] & b[7];
	assign dm_int_st0_20[12] = a[12] & b[8];
	assign dm_int_st0_21[12] = a[12] & b[9];
	assign dm_int_st0_22[12] = a[12] & b[10];
	assign dm_int_st0_23[12] = a[12] & b[11];
	assign dm_int_st0_24[12] = a[12] & b[12];
	assign dm_int_st0_25[12] = a[12] & b[13];
	assign dm_int_st0_26[12] = a[12] & b[14];
	assign dm_int_st0_27[12] = a[12] & b[15];
	assign dm_int_st0_28[12] = a[12] & b[16];
	assign dm_int_st0_29[12] = a[12] & b[17];
	assign dm_int_st0_30[12] = a[12] & b[18];
	assign dm_int_st0_31[12] = a[12] & b[19];
	assign dm_int_st0_32[11] = a[12] & b[20];
	assign dm_int_st0_33[10] = a[12] & b[21];
	assign dm_int_st0_34[9] = a[12] & b[22];
	assign dm_int_st0_35[8] = a[12] & b[23];
	assign dm_int_st0_36[7] = a[12] & b[24];
	assign dm_int_st0_37[6] = a[12] & b[25];
	assign dm_int_st0_38[5] = a[12] & b[26];
	assign dm_int_st0_39[4] = a[12] & b[27];
	assign dm_int_st0_40[3] = a[12] & b[28];
	assign dm_int_st0_41[2] = a[12] & b[29];
	assign dm_int_st0_42[1] = a[12] & b[30];
	assign dm_int_st0_43[0] = a[12] & b[31];
	assign dm_int_st0_13[13] = a[13] & b[0];
	assign dm_int_st0_14[13] = a[13] & b[1];
	assign dm_int_st0_15[13] = a[13] & b[2];
	assign dm_int_st0_16[13] = a[13] & b[3];
	assign dm_int_st0_17[13] = a[13] & b[4];
	assign dm_int_st0_18[13] = a[13] & b[5];
	assign dm_int_st0_19[13] = a[13] & b[6];
	assign dm_int_st0_20[13] = a[13] & b[7];
	assign dm_int_st0_21[13] = a[13] & b[8];
	assign dm_int_st0_22[13] = a[13] & b[9];
	assign dm_int_st0_23[13] = a[13] & b[10];
	assign dm_int_st0_24[13] = a[13] & b[11];
	assign dm_int_st0_25[13] = a[13] & b[12];
	assign dm_int_st0_26[13] = a[13] & b[13];
	assign dm_int_st0_27[13] = a[13] & b[14];
	assign dm_int_st0_28[13] = a[13] & b[15];
	assign dm_int_st0_29[13] = a[13] & b[16];
	assign dm_int_st0_30[13] = a[13] & b[17];
	assign dm_int_st0_31[13] = a[13] & b[18];
	assign dm_int_st0_32[12] = a[13] & b[19];
	assign dm_int_st0_33[11] = a[13] & b[20];
	assign dm_int_st0_34[10] = a[13] & b[21];
	assign dm_int_st0_35[9] = a[13] & b[22];
	assign dm_int_st0_36[8] = a[13] & b[23];
	assign dm_int_st0_37[7] = a[13] & b[24];
	assign dm_int_st0_38[6] = a[13] & b[25];
	assign dm_int_st0_39[5] = a[13] & b[26];
	assign dm_int_st0_40[4] = a[13] & b[27];
	assign dm_int_st0_41[3] = a[13] & b[28];
	assign dm_int_st0_42[2] = a[13] & b[29];
	assign dm_int_st0_43[1] = a[13] & b[30];
	assign dm_int_st0_44[0] = a[13] & b[31];
	assign dm_int_st0_14[14] = a[14] & b[0];
	assign dm_int_st0_15[14] = a[14] & b[1];
	assign dm_int_st0_16[14] = a[14] & b[2];
	assign dm_int_st0_17[14] = a[14] & b[3];
	assign dm_int_st0_18[14] = a[14] & b[4];
	assign dm_int_st0_19[14] = a[14] & b[5];
	assign dm_int_st0_20[14] = a[14] & b[6];
	assign dm_int_st0_21[14] = a[14] & b[7];
	assign dm_int_st0_22[14] = a[14] & b[8];
	assign dm_int_st0_23[14] = a[14] & b[9];
	assign dm_int_st0_24[14] = a[14] & b[10];
	assign dm_int_st0_25[14] = a[14] & b[11];
	assign dm_int_st0_26[14] = a[14] & b[12];
	assign dm_int_st0_27[14] = a[14] & b[13];
	assign dm_int_st0_28[14] = a[14] & b[14];
	assign dm_int_st0_29[14] = a[14] & b[15];
	assign dm_int_st0_30[14] = a[14] & b[16];
	assign dm_int_st0_31[14] = a[14] & b[17];
	assign dm_int_st0_32[13] = a[14] & b[18];
	assign dm_int_st0_33[12] = a[14] & b[19];
	assign dm_int_st0_34[11] = a[14] & b[20];
	assign dm_int_st0_35[10] = a[14] & b[21];
	assign dm_int_st0_36[9] = a[14] & b[22];
	assign dm_int_st0_37[8] = a[14] & b[23];
	assign dm_int_st0_38[7] = a[14] & b[24];
	assign dm_int_st0_39[6] = a[14] & b[25];
	assign dm_int_st0_40[5] = a[14] & b[26];
	assign dm_int_st0_41[4] = a[14] & b[27];
	assign dm_int_st0_42[3] = a[14] & b[28];
	assign dm_int_st0_43[2] = a[14] & b[29];
	assign dm_int_st0_44[1] = a[14] & b[30];
	assign dm_int_st0_45[0] = a[14] & b[31];
	assign dm_int_st0_15[15] = a[15] & b[0];
	assign dm_int_st0_16[15] = a[15] & b[1];
	assign dm_int_st0_17[15] = a[15] & b[2];
	assign dm_int_st0_18[15] = a[15] & b[3];
	assign dm_int_st0_19[15] = a[15] & b[4];
	assign dm_int_st0_20[15] = a[15] & b[5];
	assign dm_int_st0_21[15] = a[15] & b[6];
	assign dm_int_st0_22[15] = a[15] & b[7];
	assign dm_int_st0_23[15] = a[15] & b[8];
	assign dm_int_st0_24[15] = a[15] & b[9];
	assign dm_int_st0_25[15] = a[15] & b[10];
	assign dm_int_st0_26[15] = a[15] & b[11];
	assign dm_int_st0_27[15] = a[15] & b[12];
	assign dm_int_st0_28[15] = a[15] & b[13];
	assign dm_int_st0_29[15] = a[15] & b[14];
	assign dm_int_st0_30[15] = a[15] & b[15];
	assign dm_int_st0_31[15] = a[15] & b[16];
	assign dm_int_st0_32[14] = a[15] & b[17];
	assign dm_int_st0_33[13] = a[15] & b[18];
	assign dm_int_st0_34[12] = a[15] & b[19];
	assign dm_int_st0_35[11] = a[15] & b[20];
	assign dm_int_st0_36[10] = a[15] & b[21];
	assign dm_int_st0_37[9] = a[15] & b[22];
	assign dm_int_st0_38[8] = a[15] & b[23];
	assign dm_int_st0_39[7] = a[15] & b[24];
	assign dm_int_st0_40[6] = a[15] & b[25];
	assign dm_int_st0_41[5] = a[15] & b[26];
	assign dm_int_st0_42[4] = a[15] & b[27];
	assign dm_int_st0_43[3] = a[15] & b[28];
	assign dm_int_st0_44[2] = a[15] & b[29];
	assign dm_int_st0_45[1] = a[15] & b[30];
	assign dm_int_st0_46[0] = a[15] & b[31];
	assign dm_int_st0_16[16] = a[16] & b[0];
	assign dm_int_st0_17[16] = a[16] & b[1];
	assign dm_int_st0_18[16] = a[16] & b[2];
	assign dm_int_st0_19[16] = a[16] & b[3];
	assign dm_int_st0_20[16] = a[16] & b[4];
	assign dm_int_st0_21[16] = a[16] & b[5];
	assign dm_int_st0_22[16] = a[16] & b[6];
	assign dm_int_st0_23[16] = a[16] & b[7];
	assign dm_int_st0_24[16] = a[16] & b[8];
	assign dm_int_st0_25[16] = a[16] & b[9];
	assign dm_int_st0_26[16] = a[16] & b[10];
	assign dm_int_st0_27[16] = a[16] & b[11];
	assign dm_int_st0_28[16] = a[16] & b[12];
	assign dm_int_st0_29[16] = a[16] & b[13];
	assign dm_int_st0_30[16] = a[16] & b[14];
	assign dm_int_st0_31[16] = a[16] & b[15];
	assign dm_int_st0_32[15] = a[16] & b[16];
	assign dm_int_st0_33[14] = a[16] & b[17];
	assign dm_int_st0_34[13] = a[16] & b[18];
	assign dm_int_st0_35[12] = a[16] & b[19];
	assign dm_int_st0_36[11] = a[16] & b[20];
	assign dm_int_st0_37[10] = a[16] & b[21];
	assign dm_int_st0_38[9] = a[16] & b[22];
	assign dm_int_st0_39[8] = a[16] & b[23];
	assign dm_int_st0_40[7] = a[16] & b[24];
	assign dm_int_st0_41[6] = a[16] & b[25];
	assign dm_int_st0_42[5] = a[16] & b[26];
	assign dm_int_st0_43[4] = a[16] & b[27];
	assign dm_int_st0_44[3] = a[16] & b[28];
	assign dm_int_st0_45[2] = a[16] & b[29];
	assign dm_int_st0_46[1] = a[16] & b[30];
	assign dm_int_st0_47[0] = a[16] & b[31];
	assign dm_int_st0_17[17] = a[17] & b[0];
	assign dm_int_st0_18[17] = a[17] & b[1];
	assign dm_int_st0_19[17] = a[17] & b[2];
	assign dm_int_st0_20[17] = a[17] & b[3];
	assign dm_int_st0_21[17] = a[17] & b[4];
	assign dm_int_st0_22[17] = a[17] & b[5];
	assign dm_int_st0_23[17] = a[17] & b[6];
	assign dm_int_st0_24[17] = a[17] & b[7];
	assign dm_int_st0_25[17] = a[17] & b[8];
	assign dm_int_st0_26[17] = a[17] & b[9];
	assign dm_int_st0_27[17] = a[17] & b[10];
	assign dm_int_st0_28[17] = a[17] & b[11];
	assign dm_int_st0_29[17] = a[17] & b[12];
	assign dm_int_st0_30[17] = a[17] & b[13];
	assign dm_int_st0_31[17] = a[17] & b[14];
	assign dm_int_st0_32[16] = a[17] & b[15];
	assign dm_int_st0_33[15] = a[17] & b[16];
	assign dm_int_st0_34[14] = a[17] & b[17];
	assign dm_int_st0_35[13] = a[17] & b[18];
	assign dm_int_st0_36[12] = a[17] & b[19];
	assign dm_int_st0_37[11] = a[17] & b[20];
	assign dm_int_st0_38[10] = a[17] & b[21];
	assign dm_int_st0_39[9] = a[17] & b[22];
	assign dm_int_st0_40[8] = a[17] & b[23];
	assign dm_int_st0_41[7] = a[17] & b[24];
	assign dm_int_st0_42[6] = a[17] & b[25];
	assign dm_int_st0_43[5] = a[17] & b[26];
	assign dm_int_st0_44[4] = a[17] & b[27];
	assign dm_int_st0_45[3] = a[17] & b[28];
	assign dm_int_st0_46[2] = a[17] & b[29];
	assign dm_int_st0_47[1] = a[17] & b[30];
	assign dm_int_st0_48[0] = a[17] & b[31];
	assign dm_int_st0_18[18] = a[18] & b[0];
	assign dm_int_st0_19[18] = a[18] & b[1];
	assign dm_int_st0_20[18] = a[18] & b[2];
	assign dm_int_st0_21[18] = a[18] & b[3];
	assign dm_int_st0_22[18] = a[18] & b[4];
	assign dm_int_st0_23[18] = a[18] & b[5];
	assign dm_int_st0_24[18] = a[18] & b[6];
	assign dm_int_st0_25[18] = a[18] & b[7];
	assign dm_int_st0_26[18] = a[18] & b[8];
	assign dm_int_st0_27[18] = a[18] & b[9];
	assign dm_int_st0_28[18] = a[18] & b[10];
	assign dm_int_st0_29[18] = a[18] & b[11];
	assign dm_int_st0_30[18] = a[18] & b[12];
	assign dm_int_st0_31[18] = a[18] & b[13];
	assign dm_int_st0_32[17] = a[18] & b[14];
	assign dm_int_st0_33[16] = a[18] & b[15];
	assign dm_int_st0_34[15] = a[18] & b[16];
	assign dm_int_st0_35[14] = a[18] & b[17];
	assign dm_int_st0_36[13] = a[18] & b[18];
	assign dm_int_st0_37[12] = a[18] & b[19];
	assign dm_int_st0_38[11] = a[18] & b[20];
	assign dm_int_st0_39[10] = a[18] & b[21];
	assign dm_int_st0_40[9] = a[18] & b[22];
	assign dm_int_st0_41[8] = a[18] & b[23];
	assign dm_int_st0_42[7] = a[18] & b[24];
	assign dm_int_st0_43[6] = a[18] & b[25];
	assign dm_int_st0_44[5] = a[18] & b[26];
	assign dm_int_st0_45[4] = a[18] & b[27];
	assign dm_int_st0_46[3] = a[18] & b[28];
	assign dm_int_st0_47[2] = a[18] & b[29];
	assign dm_int_st0_48[1] = a[18] & b[30];
	assign dm_int_st0_49[0] = a[18] & b[31];
	assign dm_int_st0_19[19] = a[19] & b[0];
	assign dm_int_st0_20[19] = a[19] & b[1];
	assign dm_int_st0_21[19] = a[19] & b[2];
	assign dm_int_st0_22[19] = a[19] & b[3];
	assign dm_int_st0_23[19] = a[19] & b[4];
	assign dm_int_st0_24[19] = a[19] & b[5];
	assign dm_int_st0_25[19] = a[19] & b[6];
	assign dm_int_st0_26[19] = a[19] & b[7];
	assign dm_int_st0_27[19] = a[19] & b[8];
	assign dm_int_st0_28[19] = a[19] & b[9];
	assign dm_int_st0_29[19] = a[19] & b[10];
	assign dm_int_st0_30[19] = a[19] & b[11];
	assign dm_int_st0_31[19] = a[19] & b[12];
	assign dm_int_st0_32[18] = a[19] & b[13];
	assign dm_int_st0_33[17] = a[19] & b[14];
	assign dm_int_st0_34[16] = a[19] & b[15];
	assign dm_int_st0_35[15] = a[19] & b[16];
	assign dm_int_st0_36[14] = a[19] & b[17];
	assign dm_int_st0_37[13] = a[19] & b[18];
	assign dm_int_st0_38[12] = a[19] & b[19];
	assign dm_int_st0_39[11] = a[19] & b[20];
	assign dm_int_st0_40[10] = a[19] & b[21];
	assign dm_int_st0_41[9] = a[19] & b[22];
	assign dm_int_st0_42[8] = a[19] & b[23];
	assign dm_int_st0_43[7] = a[19] & b[24];
	assign dm_int_st0_44[6] = a[19] & b[25];
	assign dm_int_st0_45[5] = a[19] & b[26];
	assign dm_int_st0_46[4] = a[19] & b[27];
	assign dm_int_st0_47[3] = a[19] & b[28];
	assign dm_int_st0_48[2] = a[19] & b[29];
	assign dm_int_st0_49[1] = a[19] & b[30];
	assign dm_int_st0_50[0] = a[19] & b[31];
	assign dm_int_st0_20[20] = a[20] & b[0];
	assign dm_int_st0_21[20] = a[20] & b[1];
	assign dm_int_st0_22[20] = a[20] & b[2];
	assign dm_int_st0_23[20] = a[20] & b[3];
	assign dm_int_st0_24[20] = a[20] & b[4];
	assign dm_int_st0_25[20] = a[20] & b[5];
	assign dm_int_st0_26[20] = a[20] & b[6];
	assign dm_int_st0_27[20] = a[20] & b[7];
	assign dm_int_st0_28[20] = a[20] & b[8];
	assign dm_int_st0_29[20] = a[20] & b[9];
	assign dm_int_st0_30[20] = a[20] & b[10];
	assign dm_int_st0_31[20] = a[20] & b[11];
	assign dm_int_st0_32[19] = a[20] & b[12];
	assign dm_int_st0_33[18] = a[20] & b[13];
	assign dm_int_st0_34[17] = a[20] & b[14];
	assign dm_int_st0_35[16] = a[20] & b[15];
	assign dm_int_st0_36[15] = a[20] & b[16];
	assign dm_int_st0_37[14] = a[20] & b[17];
	assign dm_int_st0_38[13] = a[20] & b[18];
	assign dm_int_st0_39[12] = a[20] & b[19];
	assign dm_int_st0_40[11] = a[20] & b[20];
	assign dm_int_st0_41[10] = a[20] & b[21];
	assign dm_int_st0_42[9] = a[20] & b[22];
	assign dm_int_st0_43[8] = a[20] & b[23];
	assign dm_int_st0_44[7] = a[20] & b[24];
	assign dm_int_st0_45[6] = a[20] & b[25];
	assign dm_int_st0_46[5] = a[20] & b[26];
	assign dm_int_st0_47[4] = a[20] & b[27];
	assign dm_int_st0_48[3] = a[20] & b[28];
	assign dm_int_st0_49[2] = a[20] & b[29];
	assign dm_int_st0_50[1] = a[20] & b[30];
	assign dm_int_st0_51[0] = a[20] & b[31];
	assign dm_int_st0_21[21] = a[21] & b[0];
	assign dm_int_st0_22[21] = a[21] & b[1];
	assign dm_int_st0_23[21] = a[21] & b[2];
	assign dm_int_st0_24[21] = a[21] & b[3];
	assign dm_int_st0_25[21] = a[21] & b[4];
	assign dm_int_st0_26[21] = a[21] & b[5];
	assign dm_int_st0_27[21] = a[21] & b[6];
	assign dm_int_st0_28[21] = a[21] & b[7];
	assign dm_int_st0_29[21] = a[21] & b[8];
	assign dm_int_st0_30[21] = a[21] & b[9];
	assign dm_int_st0_31[21] = a[21] & b[10];
	assign dm_int_st0_32[20] = a[21] & b[11];
	assign dm_int_st0_33[19] = a[21] & b[12];
	assign dm_int_st0_34[18] = a[21] & b[13];
	assign dm_int_st0_35[17] = a[21] & b[14];
	assign dm_int_st0_36[16] = a[21] & b[15];
	assign dm_int_st0_37[15] = a[21] & b[16];
	assign dm_int_st0_38[14] = a[21] & b[17];
	assign dm_int_st0_39[13] = a[21] & b[18];
	assign dm_int_st0_40[12] = a[21] & b[19];
	assign dm_int_st0_41[11] = a[21] & b[20];
	assign dm_int_st0_42[10] = a[21] & b[21];
	assign dm_int_st0_43[9] = a[21] & b[22];
	assign dm_int_st0_44[8] = a[21] & b[23];
	assign dm_int_st0_45[7] = a[21] & b[24];
	assign dm_int_st0_46[6] = a[21] & b[25];
	assign dm_int_st0_47[5] = a[21] & b[26];
	assign dm_int_st0_48[4] = a[21] & b[27];
	assign dm_int_st0_49[3] = a[21] & b[28];
	assign dm_int_st0_50[2] = a[21] & b[29];
	assign dm_int_st0_51[1] = a[21] & b[30];
	assign dm_int_st0_52[0] = a[21] & b[31];
	assign dm_int_st0_22[22] = a[22] & b[0];
	assign dm_int_st0_23[22] = a[22] & b[1];
	assign dm_int_st0_24[22] = a[22] & b[2];
	assign dm_int_st0_25[22] = a[22] & b[3];
	assign dm_int_st0_26[22] = a[22] & b[4];
	assign dm_int_st0_27[22] = a[22] & b[5];
	assign dm_int_st0_28[22] = a[22] & b[6];
	assign dm_int_st0_29[22] = a[22] & b[7];
	assign dm_int_st0_30[22] = a[22] & b[8];
	assign dm_int_st0_31[22] = a[22] & b[9];
	assign dm_int_st0_32[21] = a[22] & b[10];
	assign dm_int_st0_33[20] = a[22] & b[11];
	assign dm_int_st0_34[19] = a[22] & b[12];
	assign dm_int_st0_35[18] = a[22] & b[13];
	assign dm_int_st0_36[17] = a[22] & b[14];
	assign dm_int_st0_37[16] = a[22] & b[15];
	assign dm_int_st0_38[15] = a[22] & b[16];
	assign dm_int_st0_39[14] = a[22] & b[17];
	assign dm_int_st0_40[13] = a[22] & b[18];
	assign dm_int_st0_41[12] = a[22] & b[19];
	assign dm_int_st0_42[11] = a[22] & b[20];
	assign dm_int_st0_43[10] = a[22] & b[21];
	assign dm_int_st0_44[9] = a[22] & b[22];
	assign dm_int_st0_45[8] = a[22] & b[23];
	assign dm_int_st0_46[7] = a[22] & b[24];
	assign dm_int_st0_47[6] = a[22] & b[25];
	assign dm_int_st0_48[5] = a[22] & b[26];
	assign dm_int_st0_49[4] = a[22] & b[27];
	assign dm_int_st0_50[3] = a[22] & b[28];
	assign dm_int_st0_51[2] = a[22] & b[29];
	assign dm_int_st0_52[1] = a[22] & b[30];
	assign dm_int_st0_53[0] = a[22] & b[31];
	assign dm_int_st0_23[23] = a[23] & b[0];
	assign dm_int_st0_24[23] = a[23] & b[1];
	assign dm_int_st0_25[23] = a[23] & b[2];
	assign dm_int_st0_26[23] = a[23] & b[3];
	assign dm_int_st0_27[23] = a[23] & b[4];
	assign dm_int_st0_28[23] = a[23] & b[5];
	assign dm_int_st0_29[23] = a[23] & b[6];
	assign dm_int_st0_30[23] = a[23] & b[7];
	assign dm_int_st0_31[23] = a[23] & b[8];
	assign dm_int_st0_32[22] = a[23] & b[9];
	assign dm_int_st0_33[21] = a[23] & b[10];
	assign dm_int_st0_34[20] = a[23] & b[11];
	assign dm_int_st0_35[19] = a[23] & b[12];
	assign dm_int_st0_36[18] = a[23] & b[13];
	assign dm_int_st0_37[17] = a[23] & b[14];
	assign dm_int_st0_38[16] = a[23] & b[15];
	assign dm_int_st0_39[15] = a[23] & b[16];
	assign dm_int_st0_40[14] = a[23] & b[17];
	assign dm_int_st0_41[13] = a[23] & b[18];
	assign dm_int_st0_42[12] = a[23] & b[19];
	assign dm_int_st0_43[11] = a[23] & b[20];
	assign dm_int_st0_44[10] = a[23] & b[21];
	assign dm_int_st0_45[9] = a[23] & b[22];
	assign dm_int_st0_46[8] = a[23] & b[23];
	assign dm_int_st0_47[7] = a[23] & b[24];
	assign dm_int_st0_48[6] = a[23] & b[25];
	assign dm_int_st0_49[5] = a[23] & b[26];
	assign dm_int_st0_50[4] = a[23] & b[27];
	assign dm_int_st0_51[3] = a[23] & b[28];
	assign dm_int_st0_52[2] = a[23] & b[29];
	assign dm_int_st0_53[1] = a[23] & b[30];
	assign dm_int_st0_54[0] = a[23] & b[31];
	assign dm_int_st0_24[24] = a[24] & b[0];
	assign dm_int_st0_25[24] = a[24] & b[1];
	assign dm_int_st0_26[24] = a[24] & b[2];
	assign dm_int_st0_27[24] = a[24] & b[3];
	assign dm_int_st0_28[24] = a[24] & b[4];
	assign dm_int_st0_29[24] = a[24] & b[5];
	assign dm_int_st0_30[24] = a[24] & b[6];
	assign dm_int_st0_31[24] = a[24] & b[7];
	assign dm_int_st0_32[23] = a[24] & b[8];
	assign dm_int_st0_33[22] = a[24] & b[9];
	assign dm_int_st0_34[21] = a[24] & b[10];
	assign dm_int_st0_35[20] = a[24] & b[11];
	assign dm_int_st0_36[19] = a[24] & b[12];
	assign dm_int_st0_37[18] = a[24] & b[13];
	assign dm_int_st0_38[17] = a[24] & b[14];
	assign dm_int_st0_39[16] = a[24] & b[15];
	assign dm_int_st0_40[15] = a[24] & b[16];
	assign dm_int_st0_41[14] = a[24] & b[17];
	assign dm_int_st0_42[13] = a[24] & b[18];
	assign dm_int_st0_43[12] = a[24] & b[19];
	assign dm_int_st0_44[11] = a[24] & b[20];
	assign dm_int_st0_45[10] = a[24] & b[21];
	assign dm_int_st0_46[9] = a[24] & b[22];
	assign dm_int_st0_47[8] = a[24] & b[23];
	assign dm_int_st0_48[7] = a[24] & b[24];
	assign dm_int_st0_49[6] = a[24] & b[25];
	assign dm_int_st0_50[5] = a[24] & b[26];
	assign dm_int_st0_51[4] = a[24] & b[27];
	assign dm_int_st0_52[3] = a[24] & b[28];
	assign dm_int_st0_53[2] = a[24] & b[29];
	assign dm_int_st0_54[1] = a[24] & b[30];
	assign dm_int_st0_55[0] = a[24] & b[31];
	assign dm_int_st0_25[25] = a[25] & b[0];
	assign dm_int_st0_26[25] = a[25] & b[1];
	assign dm_int_st0_27[25] = a[25] & b[2];
	assign dm_int_st0_28[25] = a[25] & b[3];
	assign dm_int_st0_29[25] = a[25] & b[4];
	assign dm_int_st0_30[25] = a[25] & b[5];
	assign dm_int_st0_31[25] = a[25] & b[6];
	assign dm_int_st0_32[24] = a[25] & b[7];
	assign dm_int_st0_33[23] = a[25] & b[8];
	assign dm_int_st0_34[22] = a[25] & b[9];
	assign dm_int_st0_35[21] = a[25] & b[10];
	assign dm_int_st0_36[20] = a[25] & b[11];
	assign dm_int_st0_37[19] = a[25] & b[12];
	assign dm_int_st0_38[18] = a[25] & b[13];
	assign dm_int_st0_39[17] = a[25] & b[14];
	assign dm_int_st0_40[16] = a[25] & b[15];
	assign dm_int_st0_41[15] = a[25] & b[16];
	assign dm_int_st0_42[14] = a[25] & b[17];
	assign dm_int_st0_43[13] = a[25] & b[18];
	assign dm_int_st0_44[12] = a[25] & b[19];
	assign dm_int_st0_45[11] = a[25] & b[20];
	assign dm_int_st0_46[10] = a[25] & b[21];
	assign dm_int_st0_47[9] = a[25] & b[22];
	assign dm_int_st0_48[8] = a[25] & b[23];
	assign dm_int_st0_49[7] = a[25] & b[24];
	assign dm_int_st0_50[6] = a[25] & b[25];
	assign dm_int_st0_51[5] = a[25] & b[26];
	assign dm_int_st0_52[4] = a[25] & b[27];
	assign dm_int_st0_53[3] = a[25] & b[28];
	assign dm_int_st0_54[2] = a[25] & b[29];
	assign dm_int_st0_55[1] = a[25] & b[30];
	assign dm_int_st0_56[0] = a[25] & b[31];
	assign dm_int_st0_26[26] = a[26] & b[0];
	assign dm_int_st0_27[26] = a[26] & b[1];
	assign dm_int_st0_28[26] = a[26] & b[2];
	assign dm_int_st0_29[26] = a[26] & b[3];
	assign dm_int_st0_30[26] = a[26] & b[4];
	assign dm_int_st0_31[26] = a[26] & b[5];
	assign dm_int_st0_32[25] = a[26] & b[6];
	assign dm_int_st0_33[24] = a[26] & b[7];
	assign dm_int_st0_34[23] = a[26] & b[8];
	assign dm_int_st0_35[22] = a[26] & b[9];
	assign dm_int_st0_36[21] = a[26] & b[10];
	assign dm_int_st0_37[20] = a[26] & b[11];
	assign dm_int_st0_38[19] = a[26] & b[12];
	assign dm_int_st0_39[18] = a[26] & b[13];
	assign dm_int_st0_40[17] = a[26] & b[14];
	assign dm_int_st0_41[16] = a[26] & b[15];
	assign dm_int_st0_42[15] = a[26] & b[16];
	assign dm_int_st0_43[14] = a[26] & b[17];
	assign dm_int_st0_44[13] = a[26] & b[18];
	assign dm_int_st0_45[12] = a[26] & b[19];
	assign dm_int_st0_46[11] = a[26] & b[20];
	assign dm_int_st0_47[10] = a[26] & b[21];
	assign dm_int_st0_48[9] = a[26] & b[22];
	assign dm_int_st0_49[8] = a[26] & b[23];
	assign dm_int_st0_50[7] = a[26] & b[24];
	assign dm_int_st0_51[6] = a[26] & b[25];
	assign dm_int_st0_52[5] = a[26] & b[26];
	assign dm_int_st0_53[4] = a[26] & b[27];
	assign dm_int_st0_54[3] = a[26] & b[28];
	assign dm_int_st0_55[2] = a[26] & b[29];
	assign dm_int_st0_56[1] = a[26] & b[30];
	assign dm_int_st0_57[0] = a[26] & b[31];
	assign dm_int_st0_27[27] = a[27] & b[0];
	assign dm_int_st0_28[27] = a[27] & b[1];
	assign dm_int_st0_29[27] = a[27] & b[2];
	assign dm_int_st0_30[27] = a[27] & b[3];
	assign dm_int_st0_31[27] = a[27] & b[4];
	assign dm_int_st0_32[26] = a[27] & b[5];
	assign dm_int_st0_33[25] = a[27] & b[6];
	assign dm_int_st0_34[24] = a[27] & b[7];
	assign dm_int_st0_35[23] = a[27] & b[8];
	assign dm_int_st0_36[22] = a[27] & b[9];
	assign dm_int_st0_37[21] = a[27] & b[10];
	assign dm_int_st0_38[20] = a[27] & b[11];
	assign dm_int_st0_39[19] = a[27] & b[12];
	assign dm_int_st0_40[18] = a[27] & b[13];
	assign dm_int_st0_41[17] = a[27] & b[14];
	assign dm_int_st0_42[16] = a[27] & b[15];
	assign dm_int_st0_43[15] = a[27] & b[16];
	assign dm_int_st0_44[14] = a[27] & b[17];
	assign dm_int_st0_45[13] = a[27] & b[18];
	assign dm_int_st0_46[12] = a[27] & b[19];
	assign dm_int_st0_47[11] = a[27] & b[20];
	assign dm_int_st0_48[10] = a[27] & b[21];
	assign dm_int_st0_49[9] = a[27] & b[22];
	assign dm_int_st0_50[8] = a[27] & b[23];
	assign dm_int_st0_51[7] = a[27] & b[24];
	assign dm_int_st0_52[6] = a[27] & b[25];
	assign dm_int_st0_53[5] = a[27] & b[26];
	assign dm_int_st0_54[4] = a[27] & b[27];
	assign dm_int_st0_55[3] = a[27] & b[28];
	assign dm_int_st0_56[2] = a[27] & b[29];
	assign dm_int_st0_57[1] = a[27] & b[30];
	assign dm_int_st0_58[0] = a[27] & b[31];
	assign dm_int_st0_28[28] = a[28] & b[0];
	assign dm_int_st0_29[28] = a[28] & b[1];
	assign dm_int_st0_30[28] = a[28] & b[2];
	assign dm_int_st0_31[28] = a[28] & b[3];
	assign dm_int_st0_32[27] = a[28] & b[4];
	assign dm_int_st0_33[26] = a[28] & b[5];
	assign dm_int_st0_34[25] = a[28] & b[6];
	assign dm_int_st0_35[24] = a[28] & b[7];
	assign dm_int_st0_36[23] = a[28] & b[8];
	assign dm_int_st0_37[22] = a[28] & b[9];
	assign dm_int_st0_38[21] = a[28] & b[10];
	assign dm_int_st0_39[20] = a[28] & b[11];
	assign dm_int_st0_40[19] = a[28] & b[12];
	assign dm_int_st0_41[18] = a[28] & b[13];
	assign dm_int_st0_42[17] = a[28] & b[14];
	assign dm_int_st0_43[16] = a[28] & b[15];
	assign dm_int_st0_44[15] = a[28] & b[16];
	assign dm_int_st0_45[14] = a[28] & b[17];
	assign dm_int_st0_46[13] = a[28] & b[18];
	assign dm_int_st0_47[12] = a[28] & b[19];
	assign dm_int_st0_48[11] = a[28] & b[20];
	assign dm_int_st0_49[10] = a[28] & b[21];
	assign dm_int_st0_50[9] = a[28] & b[22];
	assign dm_int_st0_51[8] = a[28] & b[23];
	assign dm_int_st0_52[7] = a[28] & b[24];
	assign dm_int_st0_53[6] = a[28] & b[25];
	assign dm_int_st0_54[5] = a[28] & b[26];
	assign dm_int_st0_55[4] = a[28] & b[27];
	assign dm_int_st0_56[3] = a[28] & b[28];
	assign dm_int_st0_57[2] = a[28] & b[29];
	assign dm_int_st0_58[1] = a[28] & b[30];
	assign dm_int_st0_59[0] = a[28] & b[31];
	assign dm_int_st0_29[29] = a[29] & b[0];
	assign dm_int_st0_30[29] = a[29] & b[1];
	assign dm_int_st0_31[29] = a[29] & b[2];
	assign dm_int_st0_32[28] = a[29] & b[3];
	assign dm_int_st0_33[27] = a[29] & b[4];
	assign dm_int_st0_34[26] = a[29] & b[5];
	assign dm_int_st0_35[25] = a[29] & b[6];
	assign dm_int_st0_36[24] = a[29] & b[7];
	assign dm_int_st0_37[23] = a[29] & b[8];
	assign dm_int_st0_38[22] = a[29] & b[9];
	assign dm_int_st0_39[21] = a[29] & b[10];
	assign dm_int_st0_40[20] = a[29] & b[11];
	assign dm_int_st0_41[19] = a[29] & b[12];
	assign dm_int_st0_42[18] = a[29] & b[13];
	assign dm_int_st0_43[17] = a[29] & b[14];
	assign dm_int_st0_44[16] = a[29] & b[15];
	assign dm_int_st0_45[15] = a[29] & b[16];
	assign dm_int_st0_46[14] = a[29] & b[17];
	assign dm_int_st0_47[13] = a[29] & b[18];
	assign dm_int_st0_48[12] = a[29] & b[19];
	assign dm_int_st0_49[11] = a[29] & b[20];
	assign dm_int_st0_50[10] = a[29] & b[21];
	assign dm_int_st0_51[9] = a[29] & b[22];
	assign dm_int_st0_52[8] = a[29] & b[23];
	assign dm_int_st0_53[7] = a[29] & b[24];
	assign dm_int_st0_54[6] = a[29] & b[25];
	assign dm_int_st0_55[5] = a[29] & b[26];
	assign dm_int_st0_56[4] = a[29] & b[27];
	assign dm_int_st0_57[3] = a[29] & b[28];
	assign dm_int_st0_58[2] = a[29] & b[29];
	assign dm_int_st0_59[1] = a[29] & b[30];
	assign dm_int_st0_60[0] = a[29] & b[31];
	assign dm_int_st0_30[30] = a[30] & b[0];
	assign dm_int_st0_31[30] = a[30] & b[1];
	assign dm_int_st0_32[29] = a[30] & b[2];
	assign dm_int_st0_33[28] = a[30] & b[3];
	assign dm_int_st0_34[27] = a[30] & b[4];
	assign dm_int_st0_35[26] = a[30] & b[5];
	assign dm_int_st0_36[25] = a[30] & b[6];
	assign dm_int_st0_37[24] = a[30] & b[7];
	assign dm_int_st0_38[23] = a[30] & b[8];
	assign dm_int_st0_39[22] = a[30] & b[9];
	assign dm_int_st0_40[21] = a[30] & b[10];
	assign dm_int_st0_41[20] = a[30] & b[11];
	assign dm_int_st0_42[19] = a[30] & b[12];
	assign dm_int_st0_43[18] = a[30] & b[13];
	assign dm_int_st0_44[17] = a[30] & b[14];
	assign dm_int_st0_45[16] = a[30] & b[15];
	assign dm_int_st0_46[15] = a[30] & b[16];
	assign dm_int_st0_47[14] = a[30] & b[17];
	assign dm_int_st0_48[13] = a[30] & b[18];
	assign dm_int_st0_49[12] = a[30] & b[19];
	assign dm_int_st0_50[11] = a[30] & b[20];
	assign dm_int_st0_51[10] = a[30] & b[21];
	assign dm_int_st0_52[9] = a[30] & b[22];
	assign dm_int_st0_53[8] = a[30] & b[23];
	assign dm_int_st0_54[7] = a[30] & b[24];
	assign dm_int_st0_55[6] = a[30] & b[25];
	assign dm_int_st0_56[5] = a[30] & b[26];
	assign dm_int_st0_57[4] = a[30] & b[27];
	assign dm_int_st0_58[3] = a[30] & b[28];
	assign dm_int_st0_59[2] = a[30] & b[29];
	assign dm_int_st0_60[1] = a[30] & b[30];
	assign dm_int_st0_61[0] = a[30] & b[31];
	assign dm_int_st0_31[31] = a[31] & b[0];
	assign dm_int_st0_32[30] = a[31] & b[1];
	assign dm_int_st0_33[29] = a[31] & b[2];
	assign dm_int_st0_34[28] = a[31] & b[3];
	assign dm_int_st0_35[27] = a[31] & b[4];
	assign dm_int_st0_36[26] = a[31] & b[5];
	assign dm_int_st0_37[25] = a[31] & b[6];
	assign dm_int_st0_38[24] = a[31] & b[7];
	assign dm_int_st0_39[23] = a[31] & b[8];
	assign dm_int_st0_40[22] = a[31] & b[9];
	assign dm_int_st0_41[21] = a[31] & b[10];
	assign dm_int_st0_42[20] = a[31] & b[11];
	assign dm_int_st0_43[19] = a[31] & b[12];
	assign dm_int_st0_44[18] = a[31] & b[13];
	assign dm_int_st0_45[17] = a[31] & b[14];
	assign dm_int_st0_46[16] = a[31] & b[15];
	assign dm_int_st0_47[15] = a[31] & b[16];
	assign dm_int_st0_48[14] = a[31] & b[17];
	assign dm_int_st0_49[13] = a[31] & b[18];
	assign dm_int_st0_50[12] = a[31] & b[19];
	assign dm_int_st0_51[11] = a[31] & b[20];
	assign dm_int_st0_52[10] = a[31] & b[21];
	assign dm_int_st0_53[9] = a[31] & b[22];
	assign dm_int_st0_54[8] = a[31] & b[23];
	assign dm_int_st0_55[7] = a[31] & b[24];
	assign dm_int_st0_56[6] = a[31] & b[25];
	assign dm_int_st0_57[5] = a[31] & b[26];
	assign dm_int_st0_58[4] = a[31] & b[27];
	assign dm_int_st0_59[3] = a[31] & b[28];
	assign dm_int_st0_60[2] = a[31] & b[29];
	assign dm_int_st0_61[1] = a[31] & b[30];
	assign dm_int_st0_62[0] = a[31] & b[31];

	//// Stage 1 ////
	wire [0:0] dm_int_st1_0;
	wire [1:0] dm_int_st1_1;
	wire [2:0] dm_int_st1_2;
	wire [3:0] dm_int_st1_3;
	wire [4:0] dm_int_st1_4;
	wire [5:0] dm_int_st1_5;
	wire [6:0] dm_int_st1_6;
	wire [7:0] dm_int_st1_7;
	wire [8:0] dm_int_st1_8;
	wire [9:0] dm_int_st1_9;
	wire [10:0] dm_int_st1_10;
	wire [11:0] dm_int_st1_11;
	wire [12:0] dm_int_st1_12;
	wire [13:0] dm_int_st1_13;
	wire [14:0] dm_int_st1_14;
	wire [15:0] dm_int_st1_15;
	wire [16:0] dm_int_st1_16;
	wire [17:0] dm_int_st1_17;
	wire [18:0] dm_int_st1_18;
	wire [19:0] dm_int_st1_19;
	wire [20:0] dm_int_st1_20;
	wire [21:0] dm_int_st1_21;
	wire [22:0] dm_int_st1_22;
	wire [23:0] dm_int_st1_23;
	wire [24:0] dm_int_st1_24;
	wire [25:0] dm_int_st1_25;
	wire [26:0] dm_int_st1_26;
	wire [27:0] dm_int_st1_27;
	wire [27:0] dm_int_st1_28;
	wire [27:0] dm_int_st1_29;
	wire [27:0] dm_int_st1_30;
	wire [27:0] dm_int_st1_31;
	wire [27:0] dm_int_st1_32;
	wire [27:0] dm_int_st1_33;
	wire [27:0] dm_int_st1_34;
	wire [27:0] dm_int_st1_35;
	wire [27:0] dm_int_st1_36;
	wire [25:0] dm_int_st1_37;
	wire [24:0] dm_int_st1_38;
	wire [23:0] dm_int_st1_39;
	wire [22:0] dm_int_st1_40;
	wire [21:0] dm_int_st1_41;
	wire [20:0] dm_int_st1_42;
	wire [19:0] dm_int_st1_43;
	wire [18:0] dm_int_st1_44;
	wire [17:0] dm_int_st1_45;
	wire [16:0] dm_int_st1_46;
	wire [15:0] dm_int_st1_47;
	wire [14:0] dm_int_st1_48;
	wire [13:0] dm_int_st1_49;
	wire [12:0] dm_int_st1_50;
	wire [11:0] dm_int_st1_51;
	wire [10:0] dm_int_st1_52;
	wire [9:0] dm_int_st1_53;
	wire [8:0] dm_int_st1_54;
	wire [7:0] dm_int_st1_55;
	wire [6:0] dm_int_st1_56;
	wire [5:0] dm_int_st1_57;
	wire [4:0] dm_int_st1_58;
	wire [3:0] dm_int_st1_59;
	wire [2:0] dm_int_st1_60;
	wire [1:0] dm_int_st1_61;
	wire [0:0] dm_int_st1_62;

	// Bit 0
	assign dm_int_st1_0[0] = dm_int_st0_0[0];
	// Bit 1
	assign dm_int_st1_1[0] = dm_int_st0_1[0];
	assign dm_int_st1_1[1] = dm_int_st0_1[1];
	// Bit 2
	assign dm_int_st1_2[0] = dm_int_st0_2[0];
	assign dm_int_st1_2[1] = dm_int_st0_2[1];
	assign dm_int_st1_2[2] = dm_int_st0_2[2];
	// Bit 3
	assign dm_int_st1_3[0] = dm_int_st0_3[0];
	assign dm_int_st1_3[1] = dm_int_st0_3[1];
	assign dm_int_st1_3[2] = dm_int_st0_3[2];
	assign dm_int_st1_3[3] = dm_int_st0_3[3];
	// Bit 4
	assign dm_int_st1_4[0] = dm_int_st0_4[0];
	assign dm_int_st1_4[1] = dm_int_st0_4[1];
	assign dm_int_st1_4[2] = dm_int_st0_4[2];
	assign dm_int_st1_4[3] = dm_int_st0_4[3];
	assign dm_int_st1_4[4] = dm_int_st0_4[4];
	// Bit 5
	assign dm_int_st1_5[0] = dm_int_st0_5[0];
	assign dm_int_st1_5[1] = dm_int_st0_5[1];
	assign dm_int_st1_5[2] = dm_int_st0_5[2];
	assign dm_int_st1_5[3] = dm_int_st0_5[3];
	assign dm_int_st1_5[4] = dm_int_st0_5[4];
	assign dm_int_st1_5[5] = dm_int_st0_5[5];
	// Bit 6
	assign dm_int_st1_6[0] = dm_int_st0_6[0];
	assign dm_int_st1_6[1] = dm_int_st0_6[1];
	assign dm_int_st1_6[2] = dm_int_st0_6[2];
	assign dm_int_st1_6[3] = dm_int_st0_6[3];
	assign dm_int_st1_6[4] = dm_int_st0_6[4];
	assign dm_int_st1_6[5] = dm_int_st0_6[5];
	assign dm_int_st1_6[6] = dm_int_st0_6[6];
	// Bit 7
	assign dm_int_st1_7[0] = dm_int_st0_7[0];
	assign dm_int_st1_7[1] = dm_int_st0_7[1];
	assign dm_int_st1_7[2] = dm_int_st0_7[2];
	assign dm_int_st1_7[3] = dm_int_st0_7[3];
	assign dm_int_st1_7[4] = dm_int_st0_7[4];
	assign dm_int_st1_7[5] = dm_int_st0_7[5];
	assign dm_int_st1_7[6] = dm_int_st0_7[6];
	assign dm_int_st1_7[7] = dm_int_st0_7[7];
	// Bit 8
	assign dm_int_st1_8[0] = dm_int_st0_8[0];
	assign dm_int_st1_8[1] = dm_int_st0_8[1];
	assign dm_int_st1_8[2] = dm_int_st0_8[2];
	assign dm_int_st1_8[3] = dm_int_st0_8[3];
	assign dm_int_st1_8[4] = dm_int_st0_8[4];
	assign dm_int_st1_8[5] = dm_int_st0_8[5];
	assign dm_int_st1_8[6] = dm_int_st0_8[6];
	assign dm_int_st1_8[7] = dm_int_st0_8[7];
	assign dm_int_st1_8[8] = dm_int_st0_8[8];
	// Bit 9
	assign dm_int_st1_9[0] = dm_int_st0_9[0];
	assign dm_int_st1_9[1] = dm_int_st0_9[1];
	assign dm_int_st1_9[2] = dm_int_st0_9[2];
	assign dm_int_st1_9[3] = dm_int_st0_9[3];
	assign dm_int_st1_9[4] = dm_int_st0_9[4];
	assign dm_int_st1_9[5] = dm_int_st0_9[5];
	assign dm_int_st1_9[6] = dm_int_st0_9[6];
	assign dm_int_st1_9[7] = dm_int_st0_9[7];
	assign dm_int_st1_9[8] = dm_int_st0_9[8];
	assign dm_int_st1_9[9] = dm_int_st0_9[9];
	// Bit 10
	assign dm_int_st1_10[0] = dm_int_st0_10[0];
	assign dm_int_st1_10[1] = dm_int_st0_10[1];
	assign dm_int_st1_10[2] = dm_int_st0_10[2];
	assign dm_int_st1_10[3] = dm_int_st0_10[3];
	assign dm_int_st1_10[4] = dm_int_st0_10[4];
	assign dm_int_st1_10[5] = dm_int_st0_10[5];
	assign dm_int_st1_10[6] = dm_int_st0_10[6];
	assign dm_int_st1_10[7] = dm_int_st0_10[7];
	assign dm_int_st1_10[8] = dm_int_st0_10[8];
	assign dm_int_st1_10[9] = dm_int_st0_10[9];
	assign dm_int_st1_10[10] = dm_int_st0_10[10];
	// Bit 11
	assign dm_int_st1_11[0] = dm_int_st0_11[0];
	assign dm_int_st1_11[1] = dm_int_st0_11[1];
	assign dm_int_st1_11[2] = dm_int_st0_11[2];
	assign dm_int_st1_11[3] = dm_int_st0_11[3];
	assign dm_int_st1_11[4] = dm_int_st0_11[4];
	assign dm_int_st1_11[5] = dm_int_st0_11[5];
	assign dm_int_st1_11[6] = dm_int_st0_11[6];
	assign dm_int_st1_11[7] = dm_int_st0_11[7];
	assign dm_int_st1_11[8] = dm_int_st0_11[8];
	assign dm_int_st1_11[9] = dm_int_st0_11[9];
	assign dm_int_st1_11[10] = dm_int_st0_11[10];
	assign dm_int_st1_11[11] = dm_int_st0_11[11];
	// Bit 12
	assign dm_int_st1_12[0] = dm_int_st0_12[0];
	assign dm_int_st1_12[1] = dm_int_st0_12[1];
	assign dm_int_st1_12[2] = dm_int_st0_12[2];
	assign dm_int_st1_12[3] = dm_int_st0_12[3];
	assign dm_int_st1_12[4] = dm_int_st0_12[4];
	assign dm_int_st1_12[5] = dm_int_st0_12[5];
	assign dm_int_st1_12[6] = dm_int_st0_12[6];
	assign dm_int_st1_12[7] = dm_int_st0_12[7];
	assign dm_int_st1_12[8] = dm_int_st0_12[8];
	assign dm_int_st1_12[9] = dm_int_st0_12[9];
	assign dm_int_st1_12[10] = dm_int_st0_12[10];
	assign dm_int_st1_12[11] = dm_int_st0_12[11];
	assign dm_int_st1_12[12] = dm_int_st0_12[12];
	// Bit 13
	assign dm_int_st1_13[0] = dm_int_st0_13[0];
	assign dm_int_st1_13[1] = dm_int_st0_13[1];
	assign dm_int_st1_13[2] = dm_int_st0_13[2];
	assign dm_int_st1_13[3] = dm_int_st0_13[3];
	assign dm_int_st1_13[4] = dm_int_st0_13[4];
	assign dm_int_st1_13[5] = dm_int_st0_13[5];
	assign dm_int_st1_13[6] = dm_int_st0_13[6];
	assign dm_int_st1_13[7] = dm_int_st0_13[7];
	assign dm_int_st1_13[8] = dm_int_st0_13[8];
	assign dm_int_st1_13[9] = dm_int_st0_13[9];
	assign dm_int_st1_13[10] = dm_int_st0_13[10];
	assign dm_int_st1_13[11] = dm_int_st0_13[11];
	assign dm_int_st1_13[12] = dm_int_st0_13[12];
	assign dm_int_st1_13[13] = dm_int_st0_13[13];
	// Bit 14
	assign dm_int_st1_14[0] = dm_int_st0_14[0];
	assign dm_int_st1_14[1] = dm_int_st0_14[1];
	assign dm_int_st1_14[2] = dm_int_st0_14[2];
	assign dm_int_st1_14[3] = dm_int_st0_14[3];
	assign dm_int_st1_14[4] = dm_int_st0_14[4];
	assign dm_int_st1_14[5] = dm_int_st0_14[5];
	assign dm_int_st1_14[6] = dm_int_st0_14[6];
	assign dm_int_st1_14[7] = dm_int_st0_14[7];
	assign dm_int_st1_14[8] = dm_int_st0_14[8];
	assign dm_int_st1_14[9] = dm_int_st0_14[9];
	assign dm_int_st1_14[10] = dm_int_st0_14[10];
	assign dm_int_st1_14[11] = dm_int_st0_14[11];
	assign dm_int_st1_14[12] = dm_int_st0_14[12];
	assign dm_int_st1_14[13] = dm_int_st0_14[13];
	assign dm_int_st1_14[14] = dm_int_st0_14[14];
	// Bit 15
	assign dm_int_st1_15[0] = dm_int_st0_15[0];
	assign dm_int_st1_15[1] = dm_int_st0_15[1];
	assign dm_int_st1_15[2] = dm_int_st0_15[2];
	assign dm_int_st1_15[3] = dm_int_st0_15[3];
	assign dm_int_st1_15[4] = dm_int_st0_15[4];
	assign dm_int_st1_15[5] = dm_int_st0_15[5];
	assign dm_int_st1_15[6] = dm_int_st0_15[6];
	assign dm_int_st1_15[7] = dm_int_st0_15[7];
	assign dm_int_st1_15[8] = dm_int_st0_15[8];
	assign dm_int_st1_15[9] = dm_int_st0_15[9];
	assign dm_int_st1_15[10] = dm_int_st0_15[10];
	assign dm_int_st1_15[11] = dm_int_st0_15[11];
	assign dm_int_st1_15[12] = dm_int_st0_15[12];
	assign dm_int_st1_15[13] = dm_int_st0_15[13];
	assign dm_int_st1_15[14] = dm_int_st0_15[14];
	assign dm_int_st1_15[15] = dm_int_st0_15[15];
	// Bit 16
	assign dm_int_st1_16[0] = dm_int_st0_16[0];
	assign dm_int_st1_16[1] = dm_int_st0_16[1];
	assign dm_int_st1_16[2] = dm_int_st0_16[2];
	assign dm_int_st1_16[3] = dm_int_st0_16[3];
	assign dm_int_st1_16[4] = dm_int_st0_16[4];
	assign dm_int_st1_16[5] = dm_int_st0_16[5];
	assign dm_int_st1_16[6] = dm_int_st0_16[6];
	assign dm_int_st1_16[7] = dm_int_st0_16[7];
	assign dm_int_st1_16[8] = dm_int_st0_16[8];
	assign dm_int_st1_16[9] = dm_int_st0_16[9];
	assign dm_int_st1_16[10] = dm_int_st0_16[10];
	assign dm_int_st1_16[11] = dm_int_st0_16[11];
	assign dm_int_st1_16[12] = dm_int_st0_16[12];
	assign dm_int_st1_16[13] = dm_int_st0_16[13];
	assign dm_int_st1_16[14] = dm_int_st0_16[14];
	assign dm_int_st1_16[15] = dm_int_st0_16[15];
	assign dm_int_st1_16[16] = dm_int_st0_16[16];
	// Bit 17
	assign dm_int_st1_17[0] = dm_int_st0_17[0];
	assign dm_int_st1_17[1] = dm_int_st0_17[1];
	assign dm_int_st1_17[2] = dm_int_st0_17[2];
	assign dm_int_st1_17[3] = dm_int_st0_17[3];
	assign dm_int_st1_17[4] = dm_int_st0_17[4];
	assign dm_int_st1_17[5] = dm_int_st0_17[5];
	assign dm_int_st1_17[6] = dm_int_st0_17[6];
	assign dm_int_st1_17[7] = dm_int_st0_17[7];
	assign dm_int_st1_17[8] = dm_int_st0_17[8];
	assign dm_int_st1_17[9] = dm_int_st0_17[9];
	assign dm_int_st1_17[10] = dm_int_st0_17[10];
	assign dm_int_st1_17[11] = dm_int_st0_17[11];
	assign dm_int_st1_17[12] = dm_int_st0_17[12];
	assign dm_int_st1_17[13] = dm_int_st0_17[13];
	assign dm_int_st1_17[14] = dm_int_st0_17[14];
	assign dm_int_st1_17[15] = dm_int_st0_17[15];
	assign dm_int_st1_17[16] = dm_int_st0_17[16];
	assign dm_int_st1_17[17] = dm_int_st0_17[17];
	// Bit 18
	assign dm_int_st1_18[0] = dm_int_st0_18[0];
	assign dm_int_st1_18[1] = dm_int_st0_18[1];
	assign dm_int_st1_18[2] = dm_int_st0_18[2];
	assign dm_int_st1_18[3] = dm_int_st0_18[3];
	assign dm_int_st1_18[4] = dm_int_st0_18[4];
	assign dm_int_st1_18[5] = dm_int_st0_18[5];
	assign dm_int_st1_18[6] = dm_int_st0_18[6];
	assign dm_int_st1_18[7] = dm_int_st0_18[7];
	assign dm_int_st1_18[8] = dm_int_st0_18[8];
	assign dm_int_st1_18[9] = dm_int_st0_18[9];
	assign dm_int_st1_18[10] = dm_int_st0_18[10];
	assign dm_int_st1_18[11] = dm_int_st0_18[11];
	assign dm_int_st1_18[12] = dm_int_st0_18[12];
	assign dm_int_st1_18[13] = dm_int_st0_18[13];
	assign dm_int_st1_18[14] = dm_int_st0_18[14];
	assign dm_int_st1_18[15] = dm_int_st0_18[15];
	assign dm_int_st1_18[16] = dm_int_st0_18[16];
	assign dm_int_st1_18[17] = dm_int_st0_18[17];
	assign dm_int_st1_18[18] = dm_int_st0_18[18];
	// Bit 19
	assign dm_int_st1_19[0] = dm_int_st0_19[0];
	assign dm_int_st1_19[1] = dm_int_st0_19[1];
	assign dm_int_st1_19[2] = dm_int_st0_19[2];
	assign dm_int_st1_19[3] = dm_int_st0_19[3];
	assign dm_int_st1_19[4] = dm_int_st0_19[4];
	assign dm_int_st1_19[5] = dm_int_st0_19[5];
	assign dm_int_st1_19[6] = dm_int_st0_19[6];
	assign dm_int_st1_19[7] = dm_int_st0_19[7];
	assign dm_int_st1_19[8] = dm_int_st0_19[8];
	assign dm_int_st1_19[9] = dm_int_st0_19[9];
	assign dm_int_st1_19[10] = dm_int_st0_19[10];
	assign dm_int_st1_19[11] = dm_int_st0_19[11];
	assign dm_int_st1_19[12] = dm_int_st0_19[12];
	assign dm_int_st1_19[13] = dm_int_st0_19[13];
	assign dm_int_st1_19[14] = dm_int_st0_19[14];
	assign dm_int_st1_19[15] = dm_int_st0_19[15];
	assign dm_int_st1_19[16] = dm_int_st0_19[16];
	assign dm_int_st1_19[17] = dm_int_st0_19[17];
	assign dm_int_st1_19[18] = dm_int_st0_19[18];
	assign dm_int_st1_19[19] = dm_int_st0_19[19];
	// Bit 20
	assign dm_int_st1_20[0] = dm_int_st0_20[0];
	assign dm_int_st1_20[1] = dm_int_st0_20[1];
	assign dm_int_st1_20[2] = dm_int_st0_20[2];
	assign dm_int_st1_20[3] = dm_int_st0_20[3];
	assign dm_int_st1_20[4] = dm_int_st0_20[4];
	assign dm_int_st1_20[5] = dm_int_st0_20[5];
	assign dm_int_st1_20[6] = dm_int_st0_20[6];
	assign dm_int_st1_20[7] = dm_int_st0_20[7];
	assign dm_int_st1_20[8] = dm_int_st0_20[8];
	assign dm_int_st1_20[9] = dm_int_st0_20[9];
	assign dm_int_st1_20[10] = dm_int_st0_20[10];
	assign dm_int_st1_20[11] = dm_int_st0_20[11];
	assign dm_int_st1_20[12] = dm_int_st0_20[12];
	assign dm_int_st1_20[13] = dm_int_st0_20[13];
	assign dm_int_st1_20[14] = dm_int_st0_20[14];
	assign dm_int_st1_20[15] = dm_int_st0_20[15];
	assign dm_int_st1_20[16] = dm_int_st0_20[16];
	assign dm_int_st1_20[17] = dm_int_st0_20[17];
	assign dm_int_st1_20[18] = dm_int_st0_20[18];
	assign dm_int_st1_20[19] = dm_int_st0_20[19];
	assign dm_int_st1_20[20] = dm_int_st0_20[20];
	// Bit 21
	assign dm_int_st1_21[0] = dm_int_st0_21[0];
	assign dm_int_st1_21[1] = dm_int_st0_21[1];
	assign dm_int_st1_21[2] = dm_int_st0_21[2];
	assign dm_int_st1_21[3] = dm_int_st0_21[3];
	assign dm_int_st1_21[4] = dm_int_st0_21[4];
	assign dm_int_st1_21[5] = dm_int_st0_21[5];
	assign dm_int_st1_21[6] = dm_int_st0_21[6];
	assign dm_int_st1_21[7] = dm_int_st0_21[7];
	assign dm_int_st1_21[8] = dm_int_st0_21[8];
	assign dm_int_st1_21[9] = dm_int_st0_21[9];
	assign dm_int_st1_21[10] = dm_int_st0_21[10];
	assign dm_int_st1_21[11] = dm_int_st0_21[11];
	assign dm_int_st1_21[12] = dm_int_st0_21[12];
	assign dm_int_st1_21[13] = dm_int_st0_21[13];
	assign dm_int_st1_21[14] = dm_int_st0_21[14];
	assign dm_int_st1_21[15] = dm_int_st0_21[15];
	assign dm_int_st1_21[16] = dm_int_st0_21[16];
	assign dm_int_st1_21[17] = dm_int_st0_21[17];
	assign dm_int_st1_21[18] = dm_int_st0_21[18];
	assign dm_int_st1_21[19] = dm_int_st0_21[19];
	assign dm_int_st1_21[20] = dm_int_st0_21[20];
	assign dm_int_st1_21[21] = dm_int_st0_21[21];
	// Bit 22
	assign dm_int_st1_22[0] = dm_int_st0_22[0];
	assign dm_int_st1_22[1] = dm_int_st0_22[1];
	assign dm_int_st1_22[2] = dm_int_st0_22[2];
	assign dm_int_st1_22[3] = dm_int_st0_22[3];
	assign dm_int_st1_22[4] = dm_int_st0_22[4];
	assign dm_int_st1_22[5] = dm_int_st0_22[5];
	assign dm_int_st1_22[6] = dm_int_st0_22[6];
	assign dm_int_st1_22[7] = dm_int_st0_22[7];
	assign dm_int_st1_22[8] = dm_int_st0_22[8];
	assign dm_int_st1_22[9] = dm_int_st0_22[9];
	assign dm_int_st1_22[10] = dm_int_st0_22[10];
	assign dm_int_st1_22[11] = dm_int_st0_22[11];
	assign dm_int_st1_22[12] = dm_int_st0_22[12];
	assign dm_int_st1_22[13] = dm_int_st0_22[13];
	assign dm_int_st1_22[14] = dm_int_st0_22[14];
	assign dm_int_st1_22[15] = dm_int_st0_22[15];
	assign dm_int_st1_22[16] = dm_int_st0_22[16];
	assign dm_int_st1_22[17] = dm_int_st0_22[17];
	assign dm_int_st1_22[18] = dm_int_st0_22[18];
	assign dm_int_st1_22[19] = dm_int_st0_22[19];
	assign dm_int_st1_22[20] = dm_int_st0_22[20];
	assign dm_int_st1_22[21] = dm_int_st0_22[21];
	assign dm_int_st1_22[22] = dm_int_st0_22[22];
	// Bit 23
	assign dm_int_st1_23[0] = dm_int_st0_23[0];
	assign dm_int_st1_23[1] = dm_int_st0_23[1];
	assign dm_int_st1_23[2] = dm_int_st0_23[2];
	assign dm_int_st1_23[3] = dm_int_st0_23[3];
	assign dm_int_st1_23[4] = dm_int_st0_23[4];
	assign dm_int_st1_23[5] = dm_int_st0_23[5];
	assign dm_int_st1_23[6] = dm_int_st0_23[6];
	assign dm_int_st1_23[7] = dm_int_st0_23[7];
	assign dm_int_st1_23[8] = dm_int_st0_23[8];
	assign dm_int_st1_23[9] = dm_int_st0_23[9];
	assign dm_int_st1_23[10] = dm_int_st0_23[10];
	assign dm_int_st1_23[11] = dm_int_st0_23[11];
	assign dm_int_st1_23[12] = dm_int_st0_23[12];
	assign dm_int_st1_23[13] = dm_int_st0_23[13];
	assign dm_int_st1_23[14] = dm_int_st0_23[14];
	assign dm_int_st1_23[15] = dm_int_st0_23[15];
	assign dm_int_st1_23[16] = dm_int_st0_23[16];
	assign dm_int_st1_23[17] = dm_int_st0_23[17];
	assign dm_int_st1_23[18] = dm_int_st0_23[18];
	assign dm_int_st1_23[19] = dm_int_st0_23[19];
	assign dm_int_st1_23[20] = dm_int_st0_23[20];
	assign dm_int_st1_23[21] = dm_int_st0_23[21];
	assign dm_int_st1_23[22] = dm_int_st0_23[22];
	assign dm_int_st1_23[23] = dm_int_st0_23[23];
	// Bit 24
	assign dm_int_st1_24[0] = dm_int_st0_24[0];
	assign dm_int_st1_24[1] = dm_int_st0_24[1];
	assign dm_int_st1_24[2] = dm_int_st0_24[2];
	assign dm_int_st1_24[3] = dm_int_st0_24[3];
	assign dm_int_st1_24[4] = dm_int_st0_24[4];
	assign dm_int_st1_24[5] = dm_int_st0_24[5];
	assign dm_int_st1_24[6] = dm_int_st0_24[6];
	assign dm_int_st1_24[7] = dm_int_st0_24[7];
	assign dm_int_st1_24[8] = dm_int_st0_24[8];
	assign dm_int_st1_24[9] = dm_int_st0_24[9];
	assign dm_int_st1_24[10] = dm_int_st0_24[10];
	assign dm_int_st1_24[11] = dm_int_st0_24[11];
	assign dm_int_st1_24[12] = dm_int_st0_24[12];
	assign dm_int_st1_24[13] = dm_int_st0_24[13];
	assign dm_int_st1_24[14] = dm_int_st0_24[14];
	assign dm_int_st1_24[15] = dm_int_st0_24[15];
	assign dm_int_st1_24[16] = dm_int_st0_24[16];
	assign dm_int_st1_24[17] = dm_int_st0_24[17];
	assign dm_int_st1_24[18] = dm_int_st0_24[18];
	assign dm_int_st1_24[19] = dm_int_st0_24[19];
	assign dm_int_st1_24[20] = dm_int_st0_24[20];
	assign dm_int_st1_24[21] = dm_int_st0_24[21];
	assign dm_int_st1_24[22] = dm_int_st0_24[22];
	assign dm_int_st1_24[23] = dm_int_st0_24[23];
	assign dm_int_st1_24[24] = dm_int_st0_24[24];
	// Bit 25
	assign dm_int_st1_25[0] = dm_int_st0_25[0];
	assign dm_int_st1_25[1] = dm_int_st0_25[1];
	assign dm_int_st1_25[2] = dm_int_st0_25[2];
	assign dm_int_st1_25[3] = dm_int_st0_25[3];
	assign dm_int_st1_25[4] = dm_int_st0_25[4];
	assign dm_int_st1_25[5] = dm_int_st0_25[5];
	assign dm_int_st1_25[6] = dm_int_st0_25[6];
	assign dm_int_st1_25[7] = dm_int_st0_25[7];
	assign dm_int_st1_25[8] = dm_int_st0_25[8];
	assign dm_int_st1_25[9] = dm_int_st0_25[9];
	assign dm_int_st1_25[10] = dm_int_st0_25[10];
	assign dm_int_st1_25[11] = dm_int_st0_25[11];
	assign dm_int_st1_25[12] = dm_int_st0_25[12];
	assign dm_int_st1_25[13] = dm_int_st0_25[13];
	assign dm_int_st1_25[14] = dm_int_st0_25[14];
	assign dm_int_st1_25[15] = dm_int_st0_25[15];
	assign dm_int_st1_25[16] = dm_int_st0_25[16];
	assign dm_int_st1_25[17] = dm_int_st0_25[17];
	assign dm_int_st1_25[18] = dm_int_st0_25[18];
	assign dm_int_st1_25[19] = dm_int_st0_25[19];
	assign dm_int_st1_25[20] = dm_int_st0_25[20];
	assign dm_int_st1_25[21] = dm_int_st0_25[21];
	assign dm_int_st1_25[22] = dm_int_st0_25[22];
	assign dm_int_st1_25[23] = dm_int_st0_25[23];
	assign dm_int_st1_25[24] = dm_int_st0_25[24];
	assign dm_int_st1_25[25] = dm_int_st0_25[25];
	// Bit 26
	assign dm_int_st1_26[0] = dm_int_st0_26[0];
	assign dm_int_st1_26[1] = dm_int_st0_26[1];
	assign dm_int_st1_26[2] = dm_int_st0_26[2];
	assign dm_int_st1_26[3] = dm_int_st0_26[3];
	assign dm_int_st1_26[4] = dm_int_st0_26[4];
	assign dm_int_st1_26[5] = dm_int_st0_26[5];
	assign dm_int_st1_26[6] = dm_int_st0_26[6];
	assign dm_int_st1_26[7] = dm_int_st0_26[7];
	assign dm_int_st1_26[8] = dm_int_st0_26[8];
	assign dm_int_st1_26[9] = dm_int_st0_26[9];
	assign dm_int_st1_26[10] = dm_int_st0_26[10];
	assign dm_int_st1_26[11] = dm_int_st0_26[11];
	assign dm_int_st1_26[12] = dm_int_st0_26[12];
	assign dm_int_st1_26[13] = dm_int_st0_26[13];
	assign dm_int_st1_26[14] = dm_int_st0_26[14];
	assign dm_int_st1_26[15] = dm_int_st0_26[15];
	assign dm_int_st1_26[16] = dm_int_st0_26[16];
	assign dm_int_st1_26[17] = dm_int_st0_26[17];
	assign dm_int_st1_26[18] = dm_int_st0_26[18];
	assign dm_int_st1_26[19] = dm_int_st0_26[19];
	assign dm_int_st1_26[20] = dm_int_st0_26[20];
	assign dm_int_st1_26[21] = dm_int_st0_26[21];
	assign dm_int_st1_26[22] = dm_int_st0_26[22];
	assign dm_int_st1_26[23] = dm_int_st0_26[23];
	assign dm_int_st1_26[24] = dm_int_st0_26[24];
	assign dm_int_st1_26[25] = dm_int_st0_26[25];
	assign dm_int_st1_26[26] = dm_int_st0_26[26];
	// Bit 27
	assign dm_int_st1_27[0] = dm_int_st0_27[0];
	assign dm_int_st1_27[1] = dm_int_st0_27[1];
	assign dm_int_st1_27[2] = dm_int_st0_27[2];
	assign dm_int_st1_27[3] = dm_int_st0_27[3];
	assign dm_int_st1_27[4] = dm_int_st0_27[4];
	assign dm_int_st1_27[5] = dm_int_st0_27[5];
	assign dm_int_st1_27[6] = dm_int_st0_27[6];
	assign dm_int_st1_27[7] = dm_int_st0_27[7];
	assign dm_int_st1_27[8] = dm_int_st0_27[8];
	assign dm_int_st1_27[9] = dm_int_st0_27[9];
	assign dm_int_st1_27[10] = dm_int_st0_27[10];
	assign dm_int_st1_27[11] = dm_int_st0_27[11];
	assign dm_int_st1_27[12] = dm_int_st0_27[12];
	assign dm_int_st1_27[13] = dm_int_st0_27[13];
	assign dm_int_st1_27[14] = dm_int_st0_27[14];
	assign dm_int_st1_27[15] = dm_int_st0_27[15];
	assign dm_int_st1_27[16] = dm_int_st0_27[16];
	assign dm_int_st1_27[17] = dm_int_st0_27[17];
	assign dm_int_st1_27[18] = dm_int_st0_27[18];
	assign dm_int_st1_27[19] = dm_int_st0_27[19];
	assign dm_int_st1_27[20] = dm_int_st0_27[20];
	assign dm_int_st1_27[21] = dm_int_st0_27[21];
	assign dm_int_st1_27[22] = dm_int_st0_27[22];
	assign dm_int_st1_27[23] = dm_int_st0_27[23];
	assign dm_int_st1_27[24] = dm_int_st0_27[24];
	assign dm_int_st1_27[25] = dm_int_st0_27[25];
	assign dm_int_st1_27[26] = dm_int_st0_27[26];
	assign dm_int_st1_27[27] = dm_int_st0_27[27];
	// Bit 28
	half_adder HA0(.a(dm_int_st0_28[0]), .b(dm_int_st0_28[1]), .s(dm_int_st1_28[0]), .cout(dm_int_st1_29[0]));
	assign dm_int_st1_28[1] = dm_int_st0_28[2];
	assign dm_int_st1_28[2] = dm_int_st0_28[3];
	assign dm_int_st1_28[3] = dm_int_st0_28[4];
	assign dm_int_st1_28[4] = dm_int_st0_28[5];
	assign dm_int_st1_28[5] = dm_int_st0_28[6];
	assign dm_int_st1_28[6] = dm_int_st0_28[7];
	assign dm_int_st1_28[7] = dm_int_st0_28[8];
	assign dm_int_st1_28[8] = dm_int_st0_28[9];
	assign dm_int_st1_28[9] = dm_int_st0_28[10];
	assign dm_int_st1_28[10] = dm_int_st0_28[11];
	assign dm_int_st1_28[11] = dm_int_st0_28[12];
	assign dm_int_st1_28[12] = dm_int_st0_28[13];
	assign dm_int_st1_28[13] = dm_int_st0_28[14];
	assign dm_int_st1_28[14] = dm_int_st0_28[15];
	assign dm_int_st1_28[15] = dm_int_st0_28[16];
	assign dm_int_st1_28[16] = dm_int_st0_28[17];
	assign dm_int_st1_28[17] = dm_int_st0_28[18];
	assign dm_int_st1_28[18] = dm_int_st0_28[19];
	assign dm_int_st1_28[19] = dm_int_st0_28[20];
	assign dm_int_st1_28[20] = dm_int_st0_28[21];
	assign dm_int_st1_28[21] = dm_int_st0_28[22];
	assign dm_int_st1_28[22] = dm_int_st0_28[23];
	assign dm_int_st1_28[23] = dm_int_st0_28[24];
	assign dm_int_st1_28[24] = dm_int_st0_28[25];
	assign dm_int_st1_28[25] = dm_int_st0_28[26];
	assign dm_int_st1_28[26] = dm_int_st0_28[27];
	assign dm_int_st1_28[27] = dm_int_st0_28[28];
	// Bit 29
	full_adder FA0(.a(dm_int_st0_29[0]), .b(dm_int_st0_29[1]), .cin(dm_int_st0_29[2]), .s(dm_int_st1_29[1]), .cout(dm_int_st1_30[0]));
	half_adder HA1(.a(dm_int_st0_29[3]), .b(dm_int_st0_29[4]), .s(dm_int_st1_29[2]), .cout(dm_int_st1_30[1]));
	assign dm_int_st1_29[3] = dm_int_st0_29[5];
	assign dm_int_st1_29[4] = dm_int_st0_29[6];
	assign dm_int_st1_29[5] = dm_int_st0_29[7];
	assign dm_int_st1_29[6] = dm_int_st0_29[8];
	assign dm_int_st1_29[7] = dm_int_st0_29[9];
	assign dm_int_st1_29[8] = dm_int_st0_29[10];
	assign dm_int_st1_29[9] = dm_int_st0_29[11];
	assign dm_int_st1_29[10] = dm_int_st0_29[12];
	assign dm_int_st1_29[11] = dm_int_st0_29[13];
	assign dm_int_st1_29[12] = dm_int_st0_29[14];
	assign dm_int_st1_29[13] = dm_int_st0_29[15];
	assign dm_int_st1_29[14] = dm_int_st0_29[16];
	assign dm_int_st1_29[15] = dm_int_st0_29[17];
	assign dm_int_st1_29[16] = dm_int_st0_29[18];
	assign dm_int_st1_29[17] = dm_int_st0_29[19];
	assign dm_int_st1_29[18] = dm_int_st0_29[20];
	assign dm_int_st1_29[19] = dm_int_st0_29[21];
	assign dm_int_st1_29[20] = dm_int_st0_29[22];
	assign dm_int_st1_29[21] = dm_int_st0_29[23];
	assign dm_int_st1_29[22] = dm_int_st0_29[24];
	assign dm_int_st1_29[23] = dm_int_st0_29[25];
	assign dm_int_st1_29[24] = dm_int_st0_29[26];
	assign dm_int_st1_29[25] = dm_int_st0_29[27];
	assign dm_int_st1_29[26] = dm_int_st0_29[28];
	assign dm_int_st1_29[27] = dm_int_st0_29[29];
	// Bit 30
	full_adder FA1(.a(dm_int_st0_30[0]), .b(dm_int_st0_30[1]), .cin(dm_int_st0_30[2]), .s(dm_int_st1_30[2]), .cout(dm_int_st1_31[0]));
	full_adder FA2(.a(dm_int_st0_30[3]), .b(dm_int_st0_30[4]), .cin(dm_int_st0_30[5]), .s(dm_int_st1_30[3]), .cout(dm_int_st1_31[1]));
	half_adder HA2(.a(dm_int_st0_30[6]), .b(dm_int_st0_30[7]), .s(dm_int_st1_30[4]), .cout(dm_int_st1_31[2]));
	assign dm_int_st1_30[5] = dm_int_st0_30[8];
	assign dm_int_st1_30[6] = dm_int_st0_30[9];
	assign dm_int_st1_30[7] = dm_int_st0_30[10];
	assign dm_int_st1_30[8] = dm_int_st0_30[11];
	assign dm_int_st1_30[9] = dm_int_st0_30[12];
	assign dm_int_st1_30[10] = dm_int_st0_30[13];
	assign dm_int_st1_30[11] = dm_int_st0_30[14];
	assign dm_int_st1_30[12] = dm_int_st0_30[15];
	assign dm_int_st1_30[13] = dm_int_st0_30[16];
	assign dm_int_st1_30[14] = dm_int_st0_30[17];
	assign dm_int_st1_30[15] = dm_int_st0_30[18];
	assign dm_int_st1_30[16] = dm_int_st0_30[19];
	assign dm_int_st1_30[17] = dm_int_st0_30[20];
	assign dm_int_st1_30[18] = dm_int_st0_30[21];
	assign dm_int_st1_30[19] = dm_int_st0_30[22];
	assign dm_int_st1_30[20] = dm_int_st0_30[23];
	assign dm_int_st1_30[21] = dm_int_st0_30[24];
	assign dm_int_st1_30[22] = dm_int_st0_30[25];
	assign dm_int_st1_30[23] = dm_int_st0_30[26];
	assign dm_int_st1_30[24] = dm_int_st0_30[27];
	assign dm_int_st1_30[25] = dm_int_st0_30[28];
	assign dm_int_st1_30[26] = dm_int_st0_30[29];
	assign dm_int_st1_30[27] = dm_int_st0_30[30];
	// Bit 31
	full_adder FA3(.a(dm_int_st0_31[0]), .b(dm_int_st0_31[1]), .cin(dm_int_st0_31[2]), .s(dm_int_st1_31[3]), .cout(dm_int_st1_32[0]));
	full_adder FA4(.a(dm_int_st0_31[3]), .b(dm_int_st0_31[4]), .cin(dm_int_st0_31[5]), .s(dm_int_st1_31[4]), .cout(dm_int_st1_32[1]));
	full_adder FA5(.a(dm_int_st0_31[6]), .b(dm_int_st0_31[7]), .cin(dm_int_st0_31[8]), .s(dm_int_st1_31[5]), .cout(dm_int_st1_32[2]));
	half_adder HA3(.a(dm_int_st0_31[9]), .b(dm_int_st0_31[10]), .s(dm_int_st1_31[6]), .cout(dm_int_st1_32[3]));
	assign dm_int_st1_31[7] = dm_int_st0_31[11];
	assign dm_int_st1_31[8] = dm_int_st0_31[12];
	assign dm_int_st1_31[9] = dm_int_st0_31[13];
	assign dm_int_st1_31[10] = dm_int_st0_31[14];
	assign dm_int_st1_31[11] = dm_int_st0_31[15];
	assign dm_int_st1_31[12] = dm_int_st0_31[16];
	assign dm_int_st1_31[13] = dm_int_st0_31[17];
	assign dm_int_st1_31[14] = dm_int_st0_31[18];
	assign dm_int_st1_31[15] = dm_int_st0_31[19];
	assign dm_int_st1_31[16] = dm_int_st0_31[20];
	assign dm_int_st1_31[17] = dm_int_st0_31[21];
	assign dm_int_st1_31[18] = dm_int_st0_31[22];
	assign dm_int_st1_31[19] = dm_int_st0_31[23];
	assign dm_int_st1_31[20] = dm_int_st0_31[24];
	assign dm_int_st1_31[21] = dm_int_st0_31[25];
	assign dm_int_st1_31[22] = dm_int_st0_31[26];
	assign dm_int_st1_31[23] = dm_int_st0_31[27];
	assign dm_int_st1_31[24] = dm_int_st0_31[28];
	assign dm_int_st1_31[25] = dm_int_st0_31[29];
	assign dm_int_st1_31[26] = dm_int_st0_31[30];
	assign dm_int_st1_31[27] = dm_int_st0_31[31];
	// Bit 32
	full_adder FA6(.a(dm_int_st0_32[0]), .b(dm_int_st0_32[1]), .cin(dm_int_st0_32[2]), .s(dm_int_st1_32[4]), .cout(dm_int_st1_33[0]));
	full_adder FA7(.a(dm_int_st0_32[3]), .b(dm_int_st0_32[4]), .cin(dm_int_st0_32[5]), .s(dm_int_st1_32[5]), .cout(dm_int_st1_33[1]));
	full_adder FA8(.a(dm_int_st0_32[6]), .b(dm_int_st0_32[7]), .cin(dm_int_st0_32[8]), .s(dm_int_st1_32[6]), .cout(dm_int_st1_33[2]));
	half_adder HA4(.a(dm_int_st0_32[9]), .b(dm_int_st0_32[10]), .s(dm_int_st1_32[7]), .cout(dm_int_st1_33[3]));
	assign dm_int_st1_32[8] = dm_int_st0_32[11];
	assign dm_int_st1_32[9] = dm_int_st0_32[12];
	assign dm_int_st1_32[10] = dm_int_st0_32[13];
	assign dm_int_st1_32[11] = dm_int_st0_32[14];
	assign dm_int_st1_32[12] = dm_int_st0_32[15];
	assign dm_int_st1_32[13] = dm_int_st0_32[16];
	assign dm_int_st1_32[14] = dm_int_st0_32[17];
	assign dm_int_st1_32[15] = dm_int_st0_32[18];
	assign dm_int_st1_32[16] = dm_int_st0_32[19];
	assign dm_int_st1_32[17] = dm_int_st0_32[20];
	assign dm_int_st1_32[18] = dm_int_st0_32[21];
	assign dm_int_st1_32[19] = dm_int_st0_32[22];
	assign dm_int_st1_32[20] = dm_int_st0_32[23];
	assign dm_int_st1_32[21] = dm_int_st0_32[24];
	assign dm_int_st1_32[22] = dm_int_st0_32[25];
	assign dm_int_st1_32[23] = dm_int_st0_32[26];
	assign dm_int_st1_32[24] = dm_int_st0_32[27];
	assign dm_int_st1_32[25] = dm_int_st0_32[28];
	assign dm_int_st1_32[26] = dm_int_st0_32[29];
	assign dm_int_st1_32[27] = dm_int_st0_32[30];
	// Bit 33
	full_adder FA9(.a(dm_int_st0_33[0]), .b(dm_int_st0_33[1]), .cin(dm_int_st0_33[2]), .s(dm_int_st1_33[4]), .cout(dm_int_st1_34[0]));
	full_adder FA10(.a(dm_int_st0_33[3]), .b(dm_int_st0_33[4]), .cin(dm_int_st0_33[5]), .s(dm_int_st1_33[5]), .cout(dm_int_st1_34[1]));
	full_adder FA11(.a(dm_int_st0_33[6]), .b(dm_int_st0_33[7]), .cin(dm_int_st0_33[8]), .s(dm_int_st1_33[6]), .cout(dm_int_st1_34[2]));
	assign dm_int_st1_33[7] = dm_int_st0_33[9];
	assign dm_int_st1_33[8] = dm_int_st0_33[10];
	assign dm_int_st1_33[9] = dm_int_st0_33[11];
	assign dm_int_st1_33[10] = dm_int_st0_33[12];
	assign dm_int_st1_33[11] = dm_int_st0_33[13];
	assign dm_int_st1_33[12] = dm_int_st0_33[14];
	assign dm_int_st1_33[13] = dm_int_st0_33[15];
	assign dm_int_st1_33[14] = dm_int_st0_33[16];
	assign dm_int_st1_33[15] = dm_int_st0_33[17];
	assign dm_int_st1_33[16] = dm_int_st0_33[18];
	assign dm_int_st1_33[17] = dm_int_st0_33[19];
	assign dm_int_st1_33[18] = dm_int_st0_33[20];
	assign dm_int_st1_33[19] = dm_int_st0_33[21];
	assign dm_int_st1_33[20] = dm_int_st0_33[22];
	assign dm_int_st1_33[21] = dm_int_st0_33[23];
	assign dm_int_st1_33[22] = dm_int_st0_33[24];
	assign dm_int_st1_33[23] = dm_int_st0_33[25];
	assign dm_int_st1_33[24] = dm_int_st0_33[26];
	assign dm_int_st1_33[25] = dm_int_st0_33[27];
	assign dm_int_st1_33[26] = dm_int_st0_33[28];
	assign dm_int_st1_33[27] = dm_int_st0_33[29];
	// Bit 34
	full_adder FA12(.a(dm_int_st0_34[0]), .b(dm_int_st0_34[1]), .cin(dm_int_st0_34[2]), .s(dm_int_st1_34[3]), .cout(dm_int_st1_35[0]));
	full_adder FA13(.a(dm_int_st0_34[3]), .b(dm_int_st0_34[4]), .cin(dm_int_st0_34[5]), .s(dm_int_st1_34[4]), .cout(dm_int_st1_35[1]));
	assign dm_int_st1_34[5] = dm_int_st0_34[6];
	assign dm_int_st1_34[6] = dm_int_st0_34[7];
	assign dm_int_st1_34[7] = dm_int_st0_34[8];
	assign dm_int_st1_34[8] = dm_int_st0_34[9];
	assign dm_int_st1_34[9] = dm_int_st0_34[10];
	assign dm_int_st1_34[10] = dm_int_st0_34[11];
	assign dm_int_st1_34[11] = dm_int_st0_34[12];
	assign dm_int_st1_34[12] = dm_int_st0_34[13];
	assign dm_int_st1_34[13] = dm_int_st0_34[14];
	assign dm_int_st1_34[14] = dm_int_st0_34[15];
	assign dm_int_st1_34[15] = dm_int_st0_34[16];
	assign dm_int_st1_34[16] = dm_int_st0_34[17];
	assign dm_int_st1_34[17] = dm_int_st0_34[18];
	assign dm_int_st1_34[18] = dm_int_st0_34[19];
	assign dm_int_st1_34[19] = dm_int_st0_34[20];
	assign dm_int_st1_34[20] = dm_int_st0_34[21];
	assign dm_int_st1_34[21] = dm_int_st0_34[22];
	assign dm_int_st1_34[22] = dm_int_st0_34[23];
	assign dm_int_st1_34[23] = dm_int_st0_34[24];
	assign dm_int_st1_34[24] = dm_int_st0_34[25];
	assign dm_int_st1_34[25] = dm_int_st0_34[26];
	assign dm_int_st1_34[26] = dm_int_st0_34[27];
	assign dm_int_st1_34[27] = dm_int_st0_34[28];
	// Bit 35
	full_adder FA14(.a(dm_int_st0_35[0]), .b(dm_int_st0_35[1]), .cin(dm_int_st0_35[2]), .s(dm_int_st1_35[2]), .cout(dm_int_st1_36[0]));
	assign dm_int_st1_35[3] = dm_int_st0_35[3];
	assign dm_int_st1_35[4] = dm_int_st0_35[4];
	assign dm_int_st1_35[5] = dm_int_st0_35[5];
	assign dm_int_st1_35[6] = dm_int_st0_35[6];
	assign dm_int_st1_35[7] = dm_int_st0_35[7];
	assign dm_int_st1_35[8] = dm_int_st0_35[8];
	assign dm_int_st1_35[9] = dm_int_st0_35[9];
	assign dm_int_st1_35[10] = dm_int_st0_35[10];
	assign dm_int_st1_35[11] = dm_int_st0_35[11];
	assign dm_int_st1_35[12] = dm_int_st0_35[12];
	assign dm_int_st1_35[13] = dm_int_st0_35[13];
	assign dm_int_st1_35[14] = dm_int_st0_35[14];
	assign dm_int_st1_35[15] = dm_int_st0_35[15];
	assign dm_int_st1_35[16] = dm_int_st0_35[16];
	assign dm_int_st1_35[17] = dm_int_st0_35[17];
	assign dm_int_st1_35[18] = dm_int_st0_35[18];
	assign dm_int_st1_35[19] = dm_int_st0_35[19];
	assign dm_int_st1_35[20] = dm_int_st0_35[20];
	assign dm_int_st1_35[21] = dm_int_st0_35[21];
	assign dm_int_st1_35[22] = dm_int_st0_35[22];
	assign dm_int_st1_35[23] = dm_int_st0_35[23];
	assign dm_int_st1_35[24] = dm_int_st0_35[24];
	assign dm_int_st1_35[25] = dm_int_st0_35[25];
	assign dm_int_st1_35[26] = dm_int_st0_35[26];
	assign dm_int_st1_35[27] = dm_int_st0_35[27];
	// Bit 36
	assign dm_int_st1_36[1] = dm_int_st0_36[0];
	assign dm_int_st1_36[2] = dm_int_st0_36[1];
	assign dm_int_st1_36[3] = dm_int_st0_36[2];
	assign dm_int_st1_36[4] = dm_int_st0_36[3];
	assign dm_int_st1_36[5] = dm_int_st0_36[4];
	assign dm_int_st1_36[6] = dm_int_st0_36[5];
	assign dm_int_st1_36[7] = dm_int_st0_36[6];
	assign dm_int_st1_36[8] = dm_int_st0_36[7];
	assign dm_int_st1_36[9] = dm_int_st0_36[8];
	assign dm_int_st1_36[10] = dm_int_st0_36[9];
	assign dm_int_st1_36[11] = dm_int_st0_36[10];
	assign dm_int_st1_36[12] = dm_int_st0_36[11];
	assign dm_int_st1_36[13] = dm_int_st0_36[12];
	assign dm_int_st1_36[14] = dm_int_st0_36[13];
	assign dm_int_st1_36[15] = dm_int_st0_36[14];
	assign dm_int_st1_36[16] = dm_int_st0_36[15];
	assign dm_int_st1_36[17] = dm_int_st0_36[16];
	assign dm_int_st1_36[18] = dm_int_st0_36[17];
	assign dm_int_st1_36[19] = dm_int_st0_36[18];
	assign dm_int_st1_36[20] = dm_int_st0_36[19];
	assign dm_int_st1_36[21] = dm_int_st0_36[20];
	assign dm_int_st1_36[22] = dm_int_st0_36[21];
	assign dm_int_st1_36[23] = dm_int_st0_36[22];
	assign dm_int_st1_36[24] = dm_int_st0_36[23];
	assign dm_int_st1_36[25] = dm_int_st0_36[24];
	assign dm_int_st1_36[26] = dm_int_st0_36[25];
	assign dm_int_st1_36[27] = dm_int_st0_36[26];
	// Bit 37
	assign dm_int_st1_37[0] = dm_int_st0_37[0];
	assign dm_int_st1_37[1] = dm_int_st0_37[1];
	assign dm_int_st1_37[2] = dm_int_st0_37[2];
	assign dm_int_st1_37[3] = dm_int_st0_37[3];
	assign dm_int_st1_37[4] = dm_int_st0_37[4];
	assign dm_int_st1_37[5] = dm_int_st0_37[5];
	assign dm_int_st1_37[6] = dm_int_st0_37[6];
	assign dm_int_st1_37[7] = dm_int_st0_37[7];
	assign dm_int_st1_37[8] = dm_int_st0_37[8];
	assign dm_int_st1_37[9] = dm_int_st0_37[9];
	assign dm_int_st1_37[10] = dm_int_st0_37[10];
	assign dm_int_st1_37[11] = dm_int_st0_37[11];
	assign dm_int_st1_37[12] = dm_int_st0_37[12];
	assign dm_int_st1_37[13] = dm_int_st0_37[13];
	assign dm_int_st1_37[14] = dm_int_st0_37[14];
	assign dm_int_st1_37[15] = dm_int_st0_37[15];
	assign dm_int_st1_37[16] = dm_int_st0_37[16];
	assign dm_int_st1_37[17] = dm_int_st0_37[17];
	assign dm_int_st1_37[18] = dm_int_st0_37[18];
	assign dm_int_st1_37[19] = dm_int_st0_37[19];
	assign dm_int_st1_37[20] = dm_int_st0_37[20];
	assign dm_int_st1_37[21] = dm_int_st0_37[21];
	assign dm_int_st1_37[22] = dm_int_st0_37[22];
	assign dm_int_st1_37[23] = dm_int_st0_37[23];
	assign dm_int_st1_37[24] = dm_int_st0_37[24];
	assign dm_int_st1_37[25] = dm_int_st0_37[25];
	// Bit 38
	assign dm_int_st1_38[0] = dm_int_st0_38[0];
	assign dm_int_st1_38[1] = dm_int_st0_38[1];
	assign dm_int_st1_38[2] = dm_int_st0_38[2];
	assign dm_int_st1_38[3] = dm_int_st0_38[3];
	assign dm_int_st1_38[4] = dm_int_st0_38[4];
	assign dm_int_st1_38[5] = dm_int_st0_38[5];
	assign dm_int_st1_38[6] = dm_int_st0_38[6];
	assign dm_int_st1_38[7] = dm_int_st0_38[7];
	assign dm_int_st1_38[8] = dm_int_st0_38[8];
	assign dm_int_st1_38[9] = dm_int_st0_38[9];
	assign dm_int_st1_38[10] = dm_int_st0_38[10];
	assign dm_int_st1_38[11] = dm_int_st0_38[11];
	assign dm_int_st1_38[12] = dm_int_st0_38[12];
	assign dm_int_st1_38[13] = dm_int_st0_38[13];
	assign dm_int_st1_38[14] = dm_int_st0_38[14];
	assign dm_int_st1_38[15] = dm_int_st0_38[15];
	assign dm_int_st1_38[16] = dm_int_st0_38[16];
	assign dm_int_st1_38[17] = dm_int_st0_38[17];
	assign dm_int_st1_38[18] = dm_int_st0_38[18];
	assign dm_int_st1_38[19] = dm_int_st0_38[19];
	assign dm_int_st1_38[20] = dm_int_st0_38[20];
	assign dm_int_st1_38[21] = dm_int_st0_38[21];
	assign dm_int_st1_38[22] = dm_int_st0_38[22];
	assign dm_int_st1_38[23] = dm_int_st0_38[23];
	assign dm_int_st1_38[24] = dm_int_st0_38[24];
	// Bit 39
	assign dm_int_st1_39[0] = dm_int_st0_39[0];
	assign dm_int_st1_39[1] = dm_int_st0_39[1];
	assign dm_int_st1_39[2] = dm_int_st0_39[2];
	assign dm_int_st1_39[3] = dm_int_st0_39[3];
	assign dm_int_st1_39[4] = dm_int_st0_39[4];
	assign dm_int_st1_39[5] = dm_int_st0_39[5];
	assign dm_int_st1_39[6] = dm_int_st0_39[6];
	assign dm_int_st1_39[7] = dm_int_st0_39[7];
	assign dm_int_st1_39[8] = dm_int_st0_39[8];
	assign dm_int_st1_39[9] = dm_int_st0_39[9];
	assign dm_int_st1_39[10] = dm_int_st0_39[10];
	assign dm_int_st1_39[11] = dm_int_st0_39[11];
	assign dm_int_st1_39[12] = dm_int_st0_39[12];
	assign dm_int_st1_39[13] = dm_int_st0_39[13];
	assign dm_int_st1_39[14] = dm_int_st0_39[14];
	assign dm_int_st1_39[15] = dm_int_st0_39[15];
	assign dm_int_st1_39[16] = dm_int_st0_39[16];
	assign dm_int_st1_39[17] = dm_int_st0_39[17];
	assign dm_int_st1_39[18] = dm_int_st0_39[18];
	assign dm_int_st1_39[19] = dm_int_st0_39[19];
	assign dm_int_st1_39[20] = dm_int_st0_39[20];
	assign dm_int_st1_39[21] = dm_int_st0_39[21];
	assign dm_int_st1_39[22] = dm_int_st0_39[22];
	assign dm_int_st1_39[23] = dm_int_st0_39[23];
	// Bit 40
	assign dm_int_st1_40[0] = dm_int_st0_40[0];
	assign dm_int_st1_40[1] = dm_int_st0_40[1];
	assign dm_int_st1_40[2] = dm_int_st0_40[2];
	assign dm_int_st1_40[3] = dm_int_st0_40[3];
	assign dm_int_st1_40[4] = dm_int_st0_40[4];
	assign dm_int_st1_40[5] = dm_int_st0_40[5];
	assign dm_int_st1_40[6] = dm_int_st0_40[6];
	assign dm_int_st1_40[7] = dm_int_st0_40[7];
	assign dm_int_st1_40[8] = dm_int_st0_40[8];
	assign dm_int_st1_40[9] = dm_int_st0_40[9];
	assign dm_int_st1_40[10] = dm_int_st0_40[10];
	assign dm_int_st1_40[11] = dm_int_st0_40[11];
	assign dm_int_st1_40[12] = dm_int_st0_40[12];
	assign dm_int_st1_40[13] = dm_int_st0_40[13];
	assign dm_int_st1_40[14] = dm_int_st0_40[14];
	assign dm_int_st1_40[15] = dm_int_st0_40[15];
	assign dm_int_st1_40[16] = dm_int_st0_40[16];
	assign dm_int_st1_40[17] = dm_int_st0_40[17];
	assign dm_int_st1_40[18] = dm_int_st0_40[18];
	assign dm_int_st1_40[19] = dm_int_st0_40[19];
	assign dm_int_st1_40[20] = dm_int_st0_40[20];
	assign dm_int_st1_40[21] = dm_int_st0_40[21];
	assign dm_int_st1_40[22] = dm_int_st0_40[22];
	// Bit 41
	assign dm_int_st1_41[0] = dm_int_st0_41[0];
	assign dm_int_st1_41[1] = dm_int_st0_41[1];
	assign dm_int_st1_41[2] = dm_int_st0_41[2];
	assign dm_int_st1_41[3] = dm_int_st0_41[3];
	assign dm_int_st1_41[4] = dm_int_st0_41[4];
	assign dm_int_st1_41[5] = dm_int_st0_41[5];
	assign dm_int_st1_41[6] = dm_int_st0_41[6];
	assign dm_int_st1_41[7] = dm_int_st0_41[7];
	assign dm_int_st1_41[8] = dm_int_st0_41[8];
	assign dm_int_st1_41[9] = dm_int_st0_41[9];
	assign dm_int_st1_41[10] = dm_int_st0_41[10];
	assign dm_int_st1_41[11] = dm_int_st0_41[11];
	assign dm_int_st1_41[12] = dm_int_st0_41[12];
	assign dm_int_st1_41[13] = dm_int_st0_41[13];
	assign dm_int_st1_41[14] = dm_int_st0_41[14];
	assign dm_int_st1_41[15] = dm_int_st0_41[15];
	assign dm_int_st1_41[16] = dm_int_st0_41[16];
	assign dm_int_st1_41[17] = dm_int_st0_41[17];
	assign dm_int_st1_41[18] = dm_int_st0_41[18];
	assign dm_int_st1_41[19] = dm_int_st0_41[19];
	assign dm_int_st1_41[20] = dm_int_st0_41[20];
	assign dm_int_st1_41[21] = dm_int_st0_41[21];
	// Bit 42
	assign dm_int_st1_42[0] = dm_int_st0_42[0];
	assign dm_int_st1_42[1] = dm_int_st0_42[1];
	assign dm_int_st1_42[2] = dm_int_st0_42[2];
	assign dm_int_st1_42[3] = dm_int_st0_42[3];
	assign dm_int_st1_42[4] = dm_int_st0_42[4];
	assign dm_int_st1_42[5] = dm_int_st0_42[5];
	assign dm_int_st1_42[6] = dm_int_st0_42[6];
	assign dm_int_st1_42[7] = dm_int_st0_42[7];
	assign dm_int_st1_42[8] = dm_int_st0_42[8];
	assign dm_int_st1_42[9] = dm_int_st0_42[9];
	assign dm_int_st1_42[10] = dm_int_st0_42[10];
	assign dm_int_st1_42[11] = dm_int_st0_42[11];
	assign dm_int_st1_42[12] = dm_int_st0_42[12];
	assign dm_int_st1_42[13] = dm_int_st0_42[13];
	assign dm_int_st1_42[14] = dm_int_st0_42[14];
	assign dm_int_st1_42[15] = dm_int_st0_42[15];
	assign dm_int_st1_42[16] = dm_int_st0_42[16];
	assign dm_int_st1_42[17] = dm_int_st0_42[17];
	assign dm_int_st1_42[18] = dm_int_st0_42[18];
	assign dm_int_st1_42[19] = dm_int_st0_42[19];
	assign dm_int_st1_42[20] = dm_int_st0_42[20];
	// Bit 43
	assign dm_int_st1_43[0] = dm_int_st0_43[0];
	assign dm_int_st1_43[1] = dm_int_st0_43[1];
	assign dm_int_st1_43[2] = dm_int_st0_43[2];
	assign dm_int_st1_43[3] = dm_int_st0_43[3];
	assign dm_int_st1_43[4] = dm_int_st0_43[4];
	assign dm_int_st1_43[5] = dm_int_st0_43[5];
	assign dm_int_st1_43[6] = dm_int_st0_43[6];
	assign dm_int_st1_43[7] = dm_int_st0_43[7];
	assign dm_int_st1_43[8] = dm_int_st0_43[8];
	assign dm_int_st1_43[9] = dm_int_st0_43[9];
	assign dm_int_st1_43[10] = dm_int_st0_43[10];
	assign dm_int_st1_43[11] = dm_int_st0_43[11];
	assign dm_int_st1_43[12] = dm_int_st0_43[12];
	assign dm_int_st1_43[13] = dm_int_st0_43[13];
	assign dm_int_st1_43[14] = dm_int_st0_43[14];
	assign dm_int_st1_43[15] = dm_int_st0_43[15];
	assign dm_int_st1_43[16] = dm_int_st0_43[16];
	assign dm_int_st1_43[17] = dm_int_st0_43[17];
	assign dm_int_st1_43[18] = dm_int_st0_43[18];
	assign dm_int_st1_43[19] = dm_int_st0_43[19];
	// Bit 44
	assign dm_int_st1_44[0] = dm_int_st0_44[0];
	assign dm_int_st1_44[1] = dm_int_st0_44[1];
	assign dm_int_st1_44[2] = dm_int_st0_44[2];
	assign dm_int_st1_44[3] = dm_int_st0_44[3];
	assign dm_int_st1_44[4] = dm_int_st0_44[4];
	assign dm_int_st1_44[5] = dm_int_st0_44[5];
	assign dm_int_st1_44[6] = dm_int_st0_44[6];
	assign dm_int_st1_44[7] = dm_int_st0_44[7];
	assign dm_int_st1_44[8] = dm_int_st0_44[8];
	assign dm_int_st1_44[9] = dm_int_st0_44[9];
	assign dm_int_st1_44[10] = dm_int_st0_44[10];
	assign dm_int_st1_44[11] = dm_int_st0_44[11];
	assign dm_int_st1_44[12] = dm_int_st0_44[12];
	assign dm_int_st1_44[13] = dm_int_st0_44[13];
	assign dm_int_st1_44[14] = dm_int_st0_44[14];
	assign dm_int_st1_44[15] = dm_int_st0_44[15];
	assign dm_int_st1_44[16] = dm_int_st0_44[16];
	assign dm_int_st1_44[17] = dm_int_st0_44[17];
	assign dm_int_st1_44[18] = dm_int_st0_44[18];
	// Bit 45
	assign dm_int_st1_45[0] = dm_int_st0_45[0];
	assign dm_int_st1_45[1] = dm_int_st0_45[1];
	assign dm_int_st1_45[2] = dm_int_st0_45[2];
	assign dm_int_st1_45[3] = dm_int_st0_45[3];
	assign dm_int_st1_45[4] = dm_int_st0_45[4];
	assign dm_int_st1_45[5] = dm_int_st0_45[5];
	assign dm_int_st1_45[6] = dm_int_st0_45[6];
	assign dm_int_st1_45[7] = dm_int_st0_45[7];
	assign dm_int_st1_45[8] = dm_int_st0_45[8];
	assign dm_int_st1_45[9] = dm_int_st0_45[9];
	assign dm_int_st1_45[10] = dm_int_st0_45[10];
	assign dm_int_st1_45[11] = dm_int_st0_45[11];
	assign dm_int_st1_45[12] = dm_int_st0_45[12];
	assign dm_int_st1_45[13] = dm_int_st0_45[13];
	assign dm_int_st1_45[14] = dm_int_st0_45[14];
	assign dm_int_st1_45[15] = dm_int_st0_45[15];
	assign dm_int_st1_45[16] = dm_int_st0_45[16];
	assign dm_int_st1_45[17] = dm_int_st0_45[17];
	// Bit 46
	assign dm_int_st1_46[0] = dm_int_st0_46[0];
	assign dm_int_st1_46[1] = dm_int_st0_46[1];
	assign dm_int_st1_46[2] = dm_int_st0_46[2];
	assign dm_int_st1_46[3] = dm_int_st0_46[3];
	assign dm_int_st1_46[4] = dm_int_st0_46[4];
	assign dm_int_st1_46[5] = dm_int_st0_46[5];
	assign dm_int_st1_46[6] = dm_int_st0_46[6];
	assign dm_int_st1_46[7] = dm_int_st0_46[7];
	assign dm_int_st1_46[8] = dm_int_st0_46[8];
	assign dm_int_st1_46[9] = dm_int_st0_46[9];
	assign dm_int_st1_46[10] = dm_int_st0_46[10];
	assign dm_int_st1_46[11] = dm_int_st0_46[11];
	assign dm_int_st1_46[12] = dm_int_st0_46[12];
	assign dm_int_st1_46[13] = dm_int_st0_46[13];
	assign dm_int_st1_46[14] = dm_int_st0_46[14];
	assign dm_int_st1_46[15] = dm_int_st0_46[15];
	assign dm_int_st1_46[16] = dm_int_st0_46[16];
	// Bit 47
	assign dm_int_st1_47[0] = dm_int_st0_47[0];
	assign dm_int_st1_47[1] = dm_int_st0_47[1];
	assign dm_int_st1_47[2] = dm_int_st0_47[2];
	assign dm_int_st1_47[3] = dm_int_st0_47[3];
	assign dm_int_st1_47[4] = dm_int_st0_47[4];
	assign dm_int_st1_47[5] = dm_int_st0_47[5];
	assign dm_int_st1_47[6] = dm_int_st0_47[6];
	assign dm_int_st1_47[7] = dm_int_st0_47[7];
	assign dm_int_st1_47[8] = dm_int_st0_47[8];
	assign dm_int_st1_47[9] = dm_int_st0_47[9];
	assign dm_int_st1_47[10] = dm_int_st0_47[10];
	assign dm_int_st1_47[11] = dm_int_st0_47[11];
	assign dm_int_st1_47[12] = dm_int_st0_47[12];
	assign dm_int_st1_47[13] = dm_int_st0_47[13];
	assign dm_int_st1_47[14] = dm_int_st0_47[14];
	assign dm_int_st1_47[15] = dm_int_st0_47[15];
	// Bit 48
	assign dm_int_st1_48[0] = dm_int_st0_48[0];
	assign dm_int_st1_48[1] = dm_int_st0_48[1];
	assign dm_int_st1_48[2] = dm_int_st0_48[2];
	assign dm_int_st1_48[3] = dm_int_st0_48[3];
	assign dm_int_st1_48[4] = dm_int_st0_48[4];
	assign dm_int_st1_48[5] = dm_int_st0_48[5];
	assign dm_int_st1_48[6] = dm_int_st0_48[6];
	assign dm_int_st1_48[7] = dm_int_st0_48[7];
	assign dm_int_st1_48[8] = dm_int_st0_48[8];
	assign dm_int_st1_48[9] = dm_int_st0_48[9];
	assign dm_int_st1_48[10] = dm_int_st0_48[10];
	assign dm_int_st1_48[11] = dm_int_st0_48[11];
	assign dm_int_st1_48[12] = dm_int_st0_48[12];
	assign dm_int_st1_48[13] = dm_int_st0_48[13];
	assign dm_int_st1_48[14] = dm_int_st0_48[14];
	// Bit 49
	assign dm_int_st1_49[0] = dm_int_st0_49[0];
	assign dm_int_st1_49[1] = dm_int_st0_49[1];
	assign dm_int_st1_49[2] = dm_int_st0_49[2];
	assign dm_int_st1_49[3] = dm_int_st0_49[3];
	assign dm_int_st1_49[4] = dm_int_st0_49[4];
	assign dm_int_st1_49[5] = dm_int_st0_49[5];
	assign dm_int_st1_49[6] = dm_int_st0_49[6];
	assign dm_int_st1_49[7] = dm_int_st0_49[7];
	assign dm_int_st1_49[8] = dm_int_st0_49[8];
	assign dm_int_st1_49[9] = dm_int_st0_49[9];
	assign dm_int_st1_49[10] = dm_int_st0_49[10];
	assign dm_int_st1_49[11] = dm_int_st0_49[11];
	assign dm_int_st1_49[12] = dm_int_st0_49[12];
	assign dm_int_st1_49[13] = dm_int_st0_49[13];
	// Bit 50
	assign dm_int_st1_50[0] = dm_int_st0_50[0];
	assign dm_int_st1_50[1] = dm_int_st0_50[1];
	assign dm_int_st1_50[2] = dm_int_st0_50[2];
	assign dm_int_st1_50[3] = dm_int_st0_50[3];
	assign dm_int_st1_50[4] = dm_int_st0_50[4];
	assign dm_int_st1_50[5] = dm_int_st0_50[5];
	assign dm_int_st1_50[6] = dm_int_st0_50[6];
	assign dm_int_st1_50[7] = dm_int_st0_50[7];
	assign dm_int_st1_50[8] = dm_int_st0_50[8];
	assign dm_int_st1_50[9] = dm_int_st0_50[9];
	assign dm_int_st1_50[10] = dm_int_st0_50[10];
	assign dm_int_st1_50[11] = dm_int_st0_50[11];
	assign dm_int_st1_50[12] = dm_int_st0_50[12];
	// Bit 51
	assign dm_int_st1_51[0] = dm_int_st0_51[0];
	assign dm_int_st1_51[1] = dm_int_st0_51[1];
	assign dm_int_st1_51[2] = dm_int_st0_51[2];
	assign dm_int_st1_51[3] = dm_int_st0_51[3];
	assign dm_int_st1_51[4] = dm_int_st0_51[4];
	assign dm_int_st1_51[5] = dm_int_st0_51[5];
	assign dm_int_st1_51[6] = dm_int_st0_51[6];
	assign dm_int_st1_51[7] = dm_int_st0_51[7];
	assign dm_int_st1_51[8] = dm_int_st0_51[8];
	assign dm_int_st1_51[9] = dm_int_st0_51[9];
	assign dm_int_st1_51[10] = dm_int_st0_51[10];
	assign dm_int_st1_51[11] = dm_int_st0_51[11];
	// Bit 52
	assign dm_int_st1_52[0] = dm_int_st0_52[0];
	assign dm_int_st1_52[1] = dm_int_st0_52[1];
	assign dm_int_st1_52[2] = dm_int_st0_52[2];
	assign dm_int_st1_52[3] = dm_int_st0_52[3];
	assign dm_int_st1_52[4] = dm_int_st0_52[4];
	assign dm_int_st1_52[5] = dm_int_st0_52[5];
	assign dm_int_st1_52[6] = dm_int_st0_52[6];
	assign dm_int_st1_52[7] = dm_int_st0_52[7];
	assign dm_int_st1_52[8] = dm_int_st0_52[8];
	assign dm_int_st1_52[9] = dm_int_st0_52[9];
	assign dm_int_st1_52[10] = dm_int_st0_52[10];
	// Bit 53
	assign dm_int_st1_53[0] = dm_int_st0_53[0];
	assign dm_int_st1_53[1] = dm_int_st0_53[1];
	assign dm_int_st1_53[2] = dm_int_st0_53[2];
	assign dm_int_st1_53[3] = dm_int_st0_53[3];
	assign dm_int_st1_53[4] = dm_int_st0_53[4];
	assign dm_int_st1_53[5] = dm_int_st0_53[5];
	assign dm_int_st1_53[6] = dm_int_st0_53[6];
	assign dm_int_st1_53[7] = dm_int_st0_53[7];
	assign dm_int_st1_53[8] = dm_int_st0_53[8];
	assign dm_int_st1_53[9] = dm_int_st0_53[9];
	// Bit 54
	assign dm_int_st1_54[0] = dm_int_st0_54[0];
	assign dm_int_st1_54[1] = dm_int_st0_54[1];
	assign dm_int_st1_54[2] = dm_int_st0_54[2];
	assign dm_int_st1_54[3] = dm_int_st0_54[3];
	assign dm_int_st1_54[4] = dm_int_st0_54[4];
	assign dm_int_st1_54[5] = dm_int_st0_54[5];
	assign dm_int_st1_54[6] = dm_int_st0_54[6];
	assign dm_int_st1_54[7] = dm_int_st0_54[7];
	assign dm_int_st1_54[8] = dm_int_st0_54[8];
	// Bit 55
	assign dm_int_st1_55[0] = dm_int_st0_55[0];
	assign dm_int_st1_55[1] = dm_int_st0_55[1];
	assign dm_int_st1_55[2] = dm_int_st0_55[2];
	assign dm_int_st1_55[3] = dm_int_st0_55[3];
	assign dm_int_st1_55[4] = dm_int_st0_55[4];
	assign dm_int_st1_55[5] = dm_int_st0_55[5];
	assign dm_int_st1_55[6] = dm_int_st0_55[6];
	assign dm_int_st1_55[7] = dm_int_st0_55[7];
	// Bit 56
	assign dm_int_st1_56[0] = dm_int_st0_56[0];
	assign dm_int_st1_56[1] = dm_int_st0_56[1];
	assign dm_int_st1_56[2] = dm_int_st0_56[2];
	assign dm_int_st1_56[3] = dm_int_st0_56[3];
	assign dm_int_st1_56[4] = dm_int_st0_56[4];
	assign dm_int_st1_56[5] = dm_int_st0_56[5];
	assign dm_int_st1_56[6] = dm_int_st0_56[6];
	// Bit 57
	assign dm_int_st1_57[0] = dm_int_st0_57[0];
	assign dm_int_st1_57[1] = dm_int_st0_57[1];
	assign dm_int_st1_57[2] = dm_int_st0_57[2];
	assign dm_int_st1_57[3] = dm_int_st0_57[3];
	assign dm_int_st1_57[4] = dm_int_st0_57[4];
	assign dm_int_st1_57[5] = dm_int_st0_57[5];
	// Bit 58
	assign dm_int_st1_58[0] = dm_int_st0_58[0];
	assign dm_int_st1_58[1] = dm_int_st0_58[1];
	assign dm_int_st1_58[2] = dm_int_st0_58[2];
	assign dm_int_st1_58[3] = dm_int_st0_58[3];
	assign dm_int_st1_58[4] = dm_int_st0_58[4];
	// Bit 59
	assign dm_int_st1_59[0] = dm_int_st0_59[0];
	assign dm_int_st1_59[1] = dm_int_st0_59[1];
	assign dm_int_st1_59[2] = dm_int_st0_59[2];
	assign dm_int_st1_59[3] = dm_int_st0_59[3];
	// Bit 60
	assign dm_int_st1_60[0] = dm_int_st0_60[0];
	assign dm_int_st1_60[1] = dm_int_st0_60[1];
	assign dm_int_st1_60[2] = dm_int_st0_60[2];
	// Bit 61
	assign dm_int_st1_61[0] = dm_int_st0_61[0];
	assign dm_int_st1_61[1] = dm_int_st0_61[1];
	// Bit 62
	assign dm_int_st1_62[0] = dm_int_st0_62[0];

	//// Stage 2 ////
	wire [0:0] dm_int_st2_0;
	wire [1:0] dm_int_st2_1;
	wire [2:0] dm_int_st2_2;
	wire [3:0] dm_int_st2_3;
	wire [4:0] dm_int_st2_4;
	wire [5:0] dm_int_st2_5;
	wire [6:0] dm_int_st2_6;
	wire [7:0] dm_int_st2_7;
	wire [8:0] dm_int_st2_8;
	wire [9:0] dm_int_st2_9;
	wire [10:0] dm_int_st2_10;
	wire [11:0] dm_int_st2_11;
	wire [12:0] dm_int_st2_12;
	wire [13:0] dm_int_st2_13;
	wire [14:0] dm_int_st2_14;
	wire [15:0] dm_int_st2_15;
	wire [16:0] dm_int_st2_16;
	wire [17:0] dm_int_st2_17;
	wire [18:0] dm_int_st2_18;
	wire [18:0] dm_int_st2_19;
	wire [18:0] dm_int_st2_20;
	wire [18:0] dm_int_st2_21;
	wire [18:0] dm_int_st2_22;
	wire [18:0] dm_int_st2_23;
	wire [18:0] dm_int_st2_24;
	wire [18:0] dm_int_st2_25;
	wire [18:0] dm_int_st2_26;
	wire [18:0] dm_int_st2_27;
	wire [18:0] dm_int_st2_28;
	wire [18:0] dm_int_st2_29;
	wire [18:0] dm_int_st2_30;
	wire [18:0] dm_int_st2_31;
	wire [18:0] dm_int_st2_32;
	wire [18:0] dm_int_st2_33;
	wire [18:0] dm_int_st2_34;
	wire [18:0] dm_int_st2_35;
	wire [18:0] dm_int_st2_36;
	wire [18:0] dm_int_st2_37;
	wire [18:0] dm_int_st2_38;
	wire [18:0] dm_int_st2_39;
	wire [18:0] dm_int_st2_40;
	wire [18:0] dm_int_st2_41;
	wire [18:0] dm_int_st2_42;
	wire [18:0] dm_int_st2_43;
	wire [18:0] dm_int_st2_44;
	wire [18:0] dm_int_st2_45;
	wire [16:0] dm_int_st2_46;
	wire [15:0] dm_int_st2_47;
	wire [14:0] dm_int_st2_48;
	wire [13:0] dm_int_st2_49;
	wire [12:0] dm_int_st2_50;
	wire [11:0] dm_int_st2_51;
	wire [10:0] dm_int_st2_52;
	wire [9:0] dm_int_st2_53;
	wire [8:0] dm_int_st2_54;
	wire [7:0] dm_int_st2_55;
	wire [6:0] dm_int_st2_56;
	wire [5:0] dm_int_st2_57;
	wire [4:0] dm_int_st2_58;
	wire [3:0] dm_int_st2_59;
	wire [2:0] dm_int_st2_60;
	wire [1:0] dm_int_st2_61;
	wire [0:0] dm_int_st2_62;

	// Bit 0
	assign dm_int_st2_0[0] = dm_int_st1_0[0];
	// Bit 1
	assign dm_int_st2_1[0] = dm_int_st1_1[0];
	assign dm_int_st2_1[1] = dm_int_st1_1[1];
	// Bit 2
	assign dm_int_st2_2[0] = dm_int_st1_2[0];
	assign dm_int_st2_2[1] = dm_int_st1_2[1];
	assign dm_int_st2_2[2] = dm_int_st1_2[2];
	// Bit 3
	assign dm_int_st2_3[0] = dm_int_st1_3[0];
	assign dm_int_st2_3[1] = dm_int_st1_3[1];
	assign dm_int_st2_3[2] = dm_int_st1_3[2];
	assign dm_int_st2_3[3] = dm_int_st1_3[3];
	// Bit 4
	assign dm_int_st2_4[0] = dm_int_st1_4[0];
	assign dm_int_st2_4[1] = dm_int_st1_4[1];
	assign dm_int_st2_4[2] = dm_int_st1_4[2];
	assign dm_int_st2_4[3] = dm_int_st1_4[3];
	assign dm_int_st2_4[4] = dm_int_st1_4[4];
	// Bit 5
	assign dm_int_st2_5[0] = dm_int_st1_5[0];
	assign dm_int_st2_5[1] = dm_int_st1_5[1];
	assign dm_int_st2_5[2] = dm_int_st1_5[2];
	assign dm_int_st2_5[3] = dm_int_st1_5[3];
	assign dm_int_st2_5[4] = dm_int_st1_5[4];
	assign dm_int_st2_5[5] = dm_int_st1_5[5];
	// Bit 6
	assign dm_int_st2_6[0] = dm_int_st1_6[0];
	assign dm_int_st2_6[1] = dm_int_st1_6[1];
	assign dm_int_st2_6[2] = dm_int_st1_6[2];
	assign dm_int_st2_6[3] = dm_int_st1_6[3];
	assign dm_int_st2_6[4] = dm_int_st1_6[4];
	assign dm_int_st2_6[5] = dm_int_st1_6[5];
	assign dm_int_st2_6[6] = dm_int_st1_6[6];
	// Bit 7
	assign dm_int_st2_7[0] = dm_int_st1_7[0];
	assign dm_int_st2_7[1] = dm_int_st1_7[1];
	assign dm_int_st2_7[2] = dm_int_st1_7[2];
	assign dm_int_st2_7[3] = dm_int_st1_7[3];
	assign dm_int_st2_7[4] = dm_int_st1_7[4];
	assign dm_int_st2_7[5] = dm_int_st1_7[5];
	assign dm_int_st2_7[6] = dm_int_st1_7[6];
	assign dm_int_st2_7[7] = dm_int_st1_7[7];
	// Bit 8
	assign dm_int_st2_8[0] = dm_int_st1_8[0];
	assign dm_int_st2_8[1] = dm_int_st1_8[1];
	assign dm_int_st2_8[2] = dm_int_st1_8[2];
	assign dm_int_st2_8[3] = dm_int_st1_8[3];
	assign dm_int_st2_8[4] = dm_int_st1_8[4];
	assign dm_int_st2_8[5] = dm_int_st1_8[5];
	assign dm_int_st2_8[6] = dm_int_st1_8[6];
	assign dm_int_st2_8[7] = dm_int_st1_8[7];
	assign dm_int_st2_8[8] = dm_int_st1_8[8];
	// Bit 9
	assign dm_int_st2_9[0] = dm_int_st1_9[0];
	assign dm_int_st2_9[1] = dm_int_st1_9[1];
	assign dm_int_st2_9[2] = dm_int_st1_9[2];
	assign dm_int_st2_9[3] = dm_int_st1_9[3];
	assign dm_int_st2_9[4] = dm_int_st1_9[4];
	assign dm_int_st2_9[5] = dm_int_st1_9[5];
	assign dm_int_st2_9[6] = dm_int_st1_9[6];
	assign dm_int_st2_9[7] = dm_int_st1_9[7];
	assign dm_int_st2_9[8] = dm_int_st1_9[8];
	assign dm_int_st2_9[9] = dm_int_st1_9[9];
	// Bit 10
	assign dm_int_st2_10[0] = dm_int_st1_10[0];
	assign dm_int_st2_10[1] = dm_int_st1_10[1];
	assign dm_int_st2_10[2] = dm_int_st1_10[2];
	assign dm_int_st2_10[3] = dm_int_st1_10[3];
	assign dm_int_st2_10[4] = dm_int_st1_10[4];
	assign dm_int_st2_10[5] = dm_int_st1_10[5];
	assign dm_int_st2_10[6] = dm_int_st1_10[6];
	assign dm_int_st2_10[7] = dm_int_st1_10[7];
	assign dm_int_st2_10[8] = dm_int_st1_10[8];
	assign dm_int_st2_10[9] = dm_int_st1_10[9];
	assign dm_int_st2_10[10] = dm_int_st1_10[10];
	// Bit 11
	assign dm_int_st2_11[0] = dm_int_st1_11[0];
	assign dm_int_st2_11[1] = dm_int_st1_11[1];
	assign dm_int_st2_11[2] = dm_int_st1_11[2];
	assign dm_int_st2_11[3] = dm_int_st1_11[3];
	assign dm_int_st2_11[4] = dm_int_st1_11[4];
	assign dm_int_st2_11[5] = dm_int_st1_11[5];
	assign dm_int_st2_11[6] = dm_int_st1_11[6];
	assign dm_int_st2_11[7] = dm_int_st1_11[7];
	assign dm_int_st2_11[8] = dm_int_st1_11[8];
	assign dm_int_st2_11[9] = dm_int_st1_11[9];
	assign dm_int_st2_11[10] = dm_int_st1_11[10];
	assign dm_int_st2_11[11] = dm_int_st1_11[11];
	// Bit 12
	assign dm_int_st2_12[0] = dm_int_st1_12[0];
	assign dm_int_st2_12[1] = dm_int_st1_12[1];
	assign dm_int_st2_12[2] = dm_int_st1_12[2];
	assign dm_int_st2_12[3] = dm_int_st1_12[3];
	assign dm_int_st2_12[4] = dm_int_st1_12[4];
	assign dm_int_st2_12[5] = dm_int_st1_12[5];
	assign dm_int_st2_12[6] = dm_int_st1_12[6];
	assign dm_int_st2_12[7] = dm_int_st1_12[7];
	assign dm_int_st2_12[8] = dm_int_st1_12[8];
	assign dm_int_st2_12[9] = dm_int_st1_12[9];
	assign dm_int_st2_12[10] = dm_int_st1_12[10];
	assign dm_int_st2_12[11] = dm_int_st1_12[11];
	assign dm_int_st2_12[12] = dm_int_st1_12[12];
	// Bit 13
	assign dm_int_st2_13[0] = dm_int_st1_13[0];
	assign dm_int_st2_13[1] = dm_int_st1_13[1];
	assign dm_int_st2_13[2] = dm_int_st1_13[2];
	assign dm_int_st2_13[3] = dm_int_st1_13[3];
	assign dm_int_st2_13[4] = dm_int_st1_13[4];
	assign dm_int_st2_13[5] = dm_int_st1_13[5];
	assign dm_int_st2_13[6] = dm_int_st1_13[6];
	assign dm_int_st2_13[7] = dm_int_st1_13[7];
	assign dm_int_st2_13[8] = dm_int_st1_13[8];
	assign dm_int_st2_13[9] = dm_int_st1_13[9];
	assign dm_int_st2_13[10] = dm_int_st1_13[10];
	assign dm_int_st2_13[11] = dm_int_st1_13[11];
	assign dm_int_st2_13[12] = dm_int_st1_13[12];
	assign dm_int_st2_13[13] = dm_int_st1_13[13];
	// Bit 14
	assign dm_int_st2_14[0] = dm_int_st1_14[0];
	assign dm_int_st2_14[1] = dm_int_st1_14[1];
	assign dm_int_st2_14[2] = dm_int_st1_14[2];
	assign dm_int_st2_14[3] = dm_int_st1_14[3];
	assign dm_int_st2_14[4] = dm_int_st1_14[4];
	assign dm_int_st2_14[5] = dm_int_st1_14[5];
	assign dm_int_st2_14[6] = dm_int_st1_14[6];
	assign dm_int_st2_14[7] = dm_int_st1_14[7];
	assign dm_int_st2_14[8] = dm_int_st1_14[8];
	assign dm_int_st2_14[9] = dm_int_st1_14[9];
	assign dm_int_st2_14[10] = dm_int_st1_14[10];
	assign dm_int_st2_14[11] = dm_int_st1_14[11];
	assign dm_int_st2_14[12] = dm_int_st1_14[12];
	assign dm_int_st2_14[13] = dm_int_st1_14[13];
	assign dm_int_st2_14[14] = dm_int_st1_14[14];
	// Bit 15
	assign dm_int_st2_15[0] = dm_int_st1_15[0];
	assign dm_int_st2_15[1] = dm_int_st1_15[1];
	assign dm_int_st2_15[2] = dm_int_st1_15[2];
	assign dm_int_st2_15[3] = dm_int_st1_15[3];
	assign dm_int_st2_15[4] = dm_int_st1_15[4];
	assign dm_int_st2_15[5] = dm_int_st1_15[5];
	assign dm_int_st2_15[6] = dm_int_st1_15[6];
	assign dm_int_st2_15[7] = dm_int_st1_15[7];
	assign dm_int_st2_15[8] = dm_int_st1_15[8];
	assign dm_int_st2_15[9] = dm_int_st1_15[9];
	assign dm_int_st2_15[10] = dm_int_st1_15[10];
	assign dm_int_st2_15[11] = dm_int_st1_15[11];
	assign dm_int_st2_15[12] = dm_int_st1_15[12];
	assign dm_int_st2_15[13] = dm_int_st1_15[13];
	assign dm_int_st2_15[14] = dm_int_st1_15[14];
	assign dm_int_st2_15[15] = dm_int_st1_15[15];
	// Bit 16
	assign dm_int_st2_16[0] = dm_int_st1_16[0];
	assign dm_int_st2_16[1] = dm_int_st1_16[1];
	assign dm_int_st2_16[2] = dm_int_st1_16[2];
	assign dm_int_st2_16[3] = dm_int_st1_16[3];
	assign dm_int_st2_16[4] = dm_int_st1_16[4];
	assign dm_int_st2_16[5] = dm_int_st1_16[5];
	assign dm_int_st2_16[6] = dm_int_st1_16[6];
	assign dm_int_st2_16[7] = dm_int_st1_16[7];
	assign dm_int_st2_16[8] = dm_int_st1_16[8];
	assign dm_int_st2_16[9] = dm_int_st1_16[9];
	assign dm_int_st2_16[10] = dm_int_st1_16[10];
	assign dm_int_st2_16[11] = dm_int_st1_16[11];
	assign dm_int_st2_16[12] = dm_int_st1_16[12];
	assign dm_int_st2_16[13] = dm_int_st1_16[13];
	assign dm_int_st2_16[14] = dm_int_st1_16[14];
	assign dm_int_st2_16[15] = dm_int_st1_16[15];
	assign dm_int_st2_16[16] = dm_int_st1_16[16];
	// Bit 17
	assign dm_int_st2_17[0] = dm_int_st1_17[0];
	assign dm_int_st2_17[1] = dm_int_st1_17[1];
	assign dm_int_st2_17[2] = dm_int_st1_17[2];
	assign dm_int_st2_17[3] = dm_int_st1_17[3];
	assign dm_int_st2_17[4] = dm_int_st1_17[4];
	assign dm_int_st2_17[5] = dm_int_st1_17[5];
	assign dm_int_st2_17[6] = dm_int_st1_17[6];
	assign dm_int_st2_17[7] = dm_int_st1_17[7];
	assign dm_int_st2_17[8] = dm_int_st1_17[8];
	assign dm_int_st2_17[9] = dm_int_st1_17[9];
	assign dm_int_st2_17[10] = dm_int_st1_17[10];
	assign dm_int_st2_17[11] = dm_int_st1_17[11];
	assign dm_int_st2_17[12] = dm_int_st1_17[12];
	assign dm_int_st2_17[13] = dm_int_st1_17[13];
	assign dm_int_st2_17[14] = dm_int_st1_17[14];
	assign dm_int_st2_17[15] = dm_int_st1_17[15];
	assign dm_int_st2_17[16] = dm_int_st1_17[16];
	assign dm_int_st2_17[17] = dm_int_st1_17[17];
	// Bit 18
	assign dm_int_st2_18[0] = dm_int_st1_18[0];
	assign dm_int_st2_18[1] = dm_int_st1_18[1];
	assign dm_int_st2_18[2] = dm_int_st1_18[2];
	assign dm_int_st2_18[3] = dm_int_st1_18[3];
	assign dm_int_st2_18[4] = dm_int_st1_18[4];
	assign dm_int_st2_18[5] = dm_int_st1_18[5];
	assign dm_int_st2_18[6] = dm_int_st1_18[6];
	assign dm_int_st2_18[7] = dm_int_st1_18[7];
	assign dm_int_st2_18[8] = dm_int_st1_18[8];
	assign dm_int_st2_18[9] = dm_int_st1_18[9];
	assign dm_int_st2_18[10] = dm_int_st1_18[10];
	assign dm_int_st2_18[11] = dm_int_st1_18[11];
	assign dm_int_st2_18[12] = dm_int_st1_18[12];
	assign dm_int_st2_18[13] = dm_int_st1_18[13];
	assign dm_int_st2_18[14] = dm_int_st1_18[14];
	assign dm_int_st2_18[15] = dm_int_st1_18[15];
	assign dm_int_st2_18[16] = dm_int_st1_18[16];
	assign dm_int_st2_18[17] = dm_int_st1_18[17];
	assign dm_int_st2_18[18] = dm_int_st1_18[18];
	// Bit 19
	half_adder HA5(.a(dm_int_st1_19[0]), .b(dm_int_st1_19[1]), .s(dm_int_st2_19[0]), .cout(dm_int_st2_20[0]));
	assign dm_int_st2_19[1] = dm_int_st1_19[2];
	assign dm_int_st2_19[2] = dm_int_st1_19[3];
	assign dm_int_st2_19[3] = dm_int_st1_19[4];
	assign dm_int_st2_19[4] = dm_int_st1_19[5];
	assign dm_int_st2_19[5] = dm_int_st1_19[6];
	assign dm_int_st2_19[6] = dm_int_st1_19[7];
	assign dm_int_st2_19[7] = dm_int_st1_19[8];
	assign dm_int_st2_19[8] = dm_int_st1_19[9];
	assign dm_int_st2_19[9] = dm_int_st1_19[10];
	assign dm_int_st2_19[10] = dm_int_st1_19[11];
	assign dm_int_st2_19[11] = dm_int_st1_19[12];
	assign dm_int_st2_19[12] = dm_int_st1_19[13];
	assign dm_int_st2_19[13] = dm_int_st1_19[14];
	assign dm_int_st2_19[14] = dm_int_st1_19[15];
	assign dm_int_st2_19[15] = dm_int_st1_19[16];
	assign dm_int_st2_19[16] = dm_int_st1_19[17];
	assign dm_int_st2_19[17] = dm_int_st1_19[18];
	assign dm_int_st2_19[18] = dm_int_st1_19[19];
	// Bit 20
	full_adder FA15(.a(dm_int_st1_20[0]), .b(dm_int_st1_20[1]), .cin(dm_int_st1_20[2]), .s(dm_int_st2_20[1]), .cout(dm_int_st2_21[0]));
	half_adder HA6(.a(dm_int_st1_20[3]), .b(dm_int_st1_20[4]), .s(dm_int_st2_20[2]), .cout(dm_int_st2_21[1]));
	assign dm_int_st2_20[3] = dm_int_st1_20[5];
	assign dm_int_st2_20[4] = dm_int_st1_20[6];
	assign dm_int_st2_20[5] = dm_int_st1_20[7];
	assign dm_int_st2_20[6] = dm_int_st1_20[8];
	assign dm_int_st2_20[7] = dm_int_st1_20[9];
	assign dm_int_st2_20[8] = dm_int_st1_20[10];
	assign dm_int_st2_20[9] = dm_int_st1_20[11];
	assign dm_int_st2_20[10] = dm_int_st1_20[12];
	assign dm_int_st2_20[11] = dm_int_st1_20[13];
	assign dm_int_st2_20[12] = dm_int_st1_20[14];
	assign dm_int_st2_20[13] = dm_int_st1_20[15];
	assign dm_int_st2_20[14] = dm_int_st1_20[16];
	assign dm_int_st2_20[15] = dm_int_st1_20[17];
	assign dm_int_st2_20[16] = dm_int_st1_20[18];
	assign dm_int_st2_20[17] = dm_int_st1_20[19];
	assign dm_int_st2_20[18] = dm_int_st1_20[20];
	// Bit 21
	full_adder FA16(.a(dm_int_st1_21[0]), .b(dm_int_st1_21[1]), .cin(dm_int_st1_21[2]), .s(dm_int_st2_21[2]), .cout(dm_int_st2_22[0]));
	full_adder FA17(.a(dm_int_st1_21[3]), .b(dm_int_st1_21[4]), .cin(dm_int_st1_21[5]), .s(dm_int_st2_21[3]), .cout(dm_int_st2_22[1]));
	half_adder HA7(.a(dm_int_st1_21[6]), .b(dm_int_st1_21[7]), .s(dm_int_st2_21[4]), .cout(dm_int_st2_22[2]));
	assign dm_int_st2_21[5] = dm_int_st1_21[8];
	assign dm_int_st2_21[6] = dm_int_st1_21[9];
	assign dm_int_st2_21[7] = dm_int_st1_21[10];
	assign dm_int_st2_21[8] = dm_int_st1_21[11];
	assign dm_int_st2_21[9] = dm_int_st1_21[12];
	assign dm_int_st2_21[10] = dm_int_st1_21[13];
	assign dm_int_st2_21[11] = dm_int_st1_21[14];
	assign dm_int_st2_21[12] = dm_int_st1_21[15];
	assign dm_int_st2_21[13] = dm_int_st1_21[16];
	assign dm_int_st2_21[14] = dm_int_st1_21[17];
	assign dm_int_st2_21[15] = dm_int_st1_21[18];
	assign dm_int_st2_21[16] = dm_int_st1_21[19];
	assign dm_int_st2_21[17] = dm_int_st1_21[20];
	assign dm_int_st2_21[18] = dm_int_st1_21[21];
	// Bit 22
	full_adder FA18(.a(dm_int_st1_22[0]), .b(dm_int_st1_22[1]), .cin(dm_int_st1_22[2]), .s(dm_int_st2_22[3]), .cout(dm_int_st2_23[0]));
	full_adder FA19(.a(dm_int_st1_22[3]), .b(dm_int_st1_22[4]), .cin(dm_int_st1_22[5]), .s(dm_int_st2_22[4]), .cout(dm_int_st2_23[1]));
	full_adder FA20(.a(dm_int_st1_22[6]), .b(dm_int_st1_22[7]), .cin(dm_int_st1_22[8]), .s(dm_int_st2_22[5]), .cout(dm_int_st2_23[2]));
	half_adder HA8(.a(dm_int_st1_22[9]), .b(dm_int_st1_22[10]), .s(dm_int_st2_22[6]), .cout(dm_int_st2_23[3]));
	assign dm_int_st2_22[7] = dm_int_st1_22[11];
	assign dm_int_st2_22[8] = dm_int_st1_22[12];
	assign dm_int_st2_22[9] = dm_int_st1_22[13];
	assign dm_int_st2_22[10] = dm_int_st1_22[14];
	assign dm_int_st2_22[11] = dm_int_st1_22[15];
	assign dm_int_st2_22[12] = dm_int_st1_22[16];
	assign dm_int_st2_22[13] = dm_int_st1_22[17];
	assign dm_int_st2_22[14] = dm_int_st1_22[18];
	assign dm_int_st2_22[15] = dm_int_st1_22[19];
	assign dm_int_st2_22[16] = dm_int_st1_22[20];
	assign dm_int_st2_22[17] = dm_int_st1_22[21];
	assign dm_int_st2_22[18] = dm_int_st1_22[22];
	// Bit 23
	full_adder FA21(.a(dm_int_st1_23[0]), .b(dm_int_st1_23[1]), .cin(dm_int_st1_23[2]), .s(dm_int_st2_23[4]), .cout(dm_int_st2_24[0]));
	full_adder FA22(.a(dm_int_st1_23[3]), .b(dm_int_st1_23[4]), .cin(dm_int_st1_23[5]), .s(dm_int_st2_23[5]), .cout(dm_int_st2_24[1]));
	full_adder FA23(.a(dm_int_st1_23[6]), .b(dm_int_st1_23[7]), .cin(dm_int_st1_23[8]), .s(dm_int_st2_23[6]), .cout(dm_int_st2_24[2]));
	full_adder FA24(.a(dm_int_st1_23[9]), .b(dm_int_st1_23[10]), .cin(dm_int_st1_23[11]), .s(dm_int_st2_23[7]), .cout(dm_int_st2_24[3]));
	half_adder HA9(.a(dm_int_st1_23[12]), .b(dm_int_st1_23[13]), .s(dm_int_st2_23[8]), .cout(dm_int_st2_24[4]));
	assign dm_int_st2_23[9] = dm_int_st1_23[14];
	assign dm_int_st2_23[10] = dm_int_st1_23[15];
	assign dm_int_st2_23[11] = dm_int_st1_23[16];
	assign dm_int_st2_23[12] = dm_int_st1_23[17];
	assign dm_int_st2_23[13] = dm_int_st1_23[18];
	assign dm_int_st2_23[14] = dm_int_st1_23[19];
	assign dm_int_st2_23[15] = dm_int_st1_23[20];
	assign dm_int_st2_23[16] = dm_int_st1_23[21];
	assign dm_int_st2_23[17] = dm_int_st1_23[22];
	assign dm_int_st2_23[18] = dm_int_st1_23[23];
	// Bit 24
	full_adder FA25(.a(dm_int_st1_24[0]), .b(dm_int_st1_24[1]), .cin(dm_int_st1_24[2]), .s(dm_int_st2_24[5]), .cout(dm_int_st2_25[0]));
	full_adder FA26(.a(dm_int_st1_24[3]), .b(dm_int_st1_24[4]), .cin(dm_int_st1_24[5]), .s(dm_int_st2_24[6]), .cout(dm_int_st2_25[1]));
	full_adder FA27(.a(dm_int_st1_24[6]), .b(dm_int_st1_24[7]), .cin(dm_int_st1_24[8]), .s(dm_int_st2_24[7]), .cout(dm_int_st2_25[2]));
	full_adder FA28(.a(dm_int_st1_24[9]), .b(dm_int_st1_24[10]), .cin(dm_int_st1_24[11]), .s(dm_int_st2_24[8]), .cout(dm_int_st2_25[3]));
	full_adder FA29(.a(dm_int_st1_24[12]), .b(dm_int_st1_24[13]), .cin(dm_int_st1_24[14]), .s(dm_int_st2_24[9]), .cout(dm_int_st2_25[4]));
	half_adder HA10(.a(dm_int_st1_24[15]), .b(dm_int_st1_24[16]), .s(dm_int_st2_24[10]), .cout(dm_int_st2_25[5]));
	assign dm_int_st2_24[11] = dm_int_st1_24[17];
	assign dm_int_st2_24[12] = dm_int_st1_24[18];
	assign dm_int_st2_24[13] = dm_int_st1_24[19];
	assign dm_int_st2_24[14] = dm_int_st1_24[20];
	assign dm_int_st2_24[15] = dm_int_st1_24[21];
	assign dm_int_st2_24[16] = dm_int_st1_24[22];
	assign dm_int_st2_24[17] = dm_int_st1_24[23];
	assign dm_int_st2_24[18] = dm_int_st1_24[24];
	// Bit 25
	full_adder FA30(.a(dm_int_st1_25[0]), .b(dm_int_st1_25[1]), .cin(dm_int_st1_25[2]), .s(dm_int_st2_25[6]), .cout(dm_int_st2_26[0]));
	full_adder FA31(.a(dm_int_st1_25[3]), .b(dm_int_st1_25[4]), .cin(dm_int_st1_25[5]), .s(dm_int_st2_25[7]), .cout(dm_int_st2_26[1]));
	full_adder FA32(.a(dm_int_st1_25[6]), .b(dm_int_st1_25[7]), .cin(dm_int_st1_25[8]), .s(dm_int_st2_25[8]), .cout(dm_int_st2_26[2]));
	full_adder FA33(.a(dm_int_st1_25[9]), .b(dm_int_st1_25[10]), .cin(dm_int_st1_25[11]), .s(dm_int_st2_25[9]), .cout(dm_int_st2_26[3]));
	full_adder FA34(.a(dm_int_st1_25[12]), .b(dm_int_st1_25[13]), .cin(dm_int_st1_25[14]), .s(dm_int_st2_25[10]), .cout(dm_int_st2_26[4]));
	full_adder FA35(.a(dm_int_st1_25[15]), .b(dm_int_st1_25[16]), .cin(dm_int_st1_25[17]), .s(dm_int_st2_25[11]), .cout(dm_int_st2_26[5]));
	half_adder HA11(.a(dm_int_st1_25[18]), .b(dm_int_st1_25[19]), .s(dm_int_st2_25[12]), .cout(dm_int_st2_26[6]));
	assign dm_int_st2_25[13] = dm_int_st1_25[20];
	assign dm_int_st2_25[14] = dm_int_st1_25[21];
	assign dm_int_st2_25[15] = dm_int_st1_25[22];
	assign dm_int_st2_25[16] = dm_int_st1_25[23];
	assign dm_int_st2_25[17] = dm_int_st1_25[24];
	assign dm_int_st2_25[18] = dm_int_st1_25[25];
	// Bit 26
	full_adder FA36(.a(dm_int_st1_26[0]), .b(dm_int_st1_26[1]), .cin(dm_int_st1_26[2]), .s(dm_int_st2_26[7]), .cout(dm_int_st2_27[0]));
	full_adder FA37(.a(dm_int_st1_26[3]), .b(dm_int_st1_26[4]), .cin(dm_int_st1_26[5]), .s(dm_int_st2_26[8]), .cout(dm_int_st2_27[1]));
	full_adder FA38(.a(dm_int_st1_26[6]), .b(dm_int_st1_26[7]), .cin(dm_int_st1_26[8]), .s(dm_int_st2_26[9]), .cout(dm_int_st2_27[2]));
	full_adder FA39(.a(dm_int_st1_26[9]), .b(dm_int_st1_26[10]), .cin(dm_int_st1_26[11]), .s(dm_int_st2_26[10]), .cout(dm_int_st2_27[3]));
	full_adder FA40(.a(dm_int_st1_26[12]), .b(dm_int_st1_26[13]), .cin(dm_int_st1_26[14]), .s(dm_int_st2_26[11]), .cout(dm_int_st2_27[4]));
	full_adder FA41(.a(dm_int_st1_26[15]), .b(dm_int_st1_26[16]), .cin(dm_int_st1_26[17]), .s(dm_int_st2_26[12]), .cout(dm_int_st2_27[5]));
	full_adder FA42(.a(dm_int_st1_26[18]), .b(dm_int_st1_26[19]), .cin(dm_int_st1_26[20]), .s(dm_int_st2_26[13]), .cout(dm_int_st2_27[6]));
	half_adder HA12(.a(dm_int_st1_26[21]), .b(dm_int_st1_26[22]), .s(dm_int_st2_26[14]), .cout(dm_int_st2_27[7]));
	assign dm_int_st2_26[15] = dm_int_st1_26[23];
	assign dm_int_st2_26[16] = dm_int_st1_26[24];
	assign dm_int_st2_26[17] = dm_int_st1_26[25];
	assign dm_int_st2_26[18] = dm_int_st1_26[26];
	// Bit 27
	full_adder FA43(.a(dm_int_st1_27[0]), .b(dm_int_st1_27[1]), .cin(dm_int_st1_27[2]), .s(dm_int_st2_27[8]), .cout(dm_int_st2_28[0]));
	full_adder FA44(.a(dm_int_st1_27[3]), .b(dm_int_st1_27[4]), .cin(dm_int_st1_27[5]), .s(dm_int_st2_27[9]), .cout(dm_int_st2_28[1]));
	full_adder FA45(.a(dm_int_st1_27[6]), .b(dm_int_st1_27[7]), .cin(dm_int_st1_27[8]), .s(dm_int_st2_27[10]), .cout(dm_int_st2_28[2]));
	full_adder FA46(.a(dm_int_st1_27[9]), .b(dm_int_st1_27[10]), .cin(dm_int_st1_27[11]), .s(dm_int_st2_27[11]), .cout(dm_int_st2_28[3]));
	full_adder FA47(.a(dm_int_st1_27[12]), .b(dm_int_st1_27[13]), .cin(dm_int_st1_27[14]), .s(dm_int_st2_27[12]), .cout(dm_int_st2_28[4]));
	full_adder FA48(.a(dm_int_st1_27[15]), .b(dm_int_st1_27[16]), .cin(dm_int_st1_27[17]), .s(dm_int_st2_27[13]), .cout(dm_int_st2_28[5]));
	full_adder FA49(.a(dm_int_st1_27[18]), .b(dm_int_st1_27[19]), .cin(dm_int_st1_27[20]), .s(dm_int_st2_27[14]), .cout(dm_int_st2_28[6]));
	full_adder FA50(.a(dm_int_st1_27[21]), .b(dm_int_st1_27[22]), .cin(dm_int_st1_27[23]), .s(dm_int_st2_27[15]), .cout(dm_int_st2_28[7]));
	half_adder HA13(.a(dm_int_st1_27[24]), .b(dm_int_st1_27[25]), .s(dm_int_st2_27[16]), .cout(dm_int_st2_28[8]));
	assign dm_int_st2_27[17] = dm_int_st1_27[26];
	assign dm_int_st2_27[18] = dm_int_st1_27[27];
	// Bit 28
	full_adder FA51(.a(dm_int_st1_28[0]), .b(dm_int_st1_28[1]), .cin(dm_int_st1_28[2]), .s(dm_int_st2_28[9]), .cout(dm_int_st2_29[0]));
	full_adder FA52(.a(dm_int_st1_28[3]), .b(dm_int_st1_28[4]), .cin(dm_int_st1_28[5]), .s(dm_int_st2_28[10]), .cout(dm_int_st2_29[1]));
	full_adder FA53(.a(dm_int_st1_28[6]), .b(dm_int_st1_28[7]), .cin(dm_int_st1_28[8]), .s(dm_int_st2_28[11]), .cout(dm_int_st2_29[2]));
	full_adder FA54(.a(dm_int_st1_28[9]), .b(dm_int_st1_28[10]), .cin(dm_int_st1_28[11]), .s(dm_int_st2_28[12]), .cout(dm_int_st2_29[3]));
	full_adder FA55(.a(dm_int_st1_28[12]), .b(dm_int_st1_28[13]), .cin(dm_int_st1_28[14]), .s(dm_int_st2_28[13]), .cout(dm_int_st2_29[4]));
	full_adder FA56(.a(dm_int_st1_28[15]), .b(dm_int_st1_28[16]), .cin(dm_int_st1_28[17]), .s(dm_int_st2_28[14]), .cout(dm_int_st2_29[5]));
	full_adder FA57(.a(dm_int_st1_28[18]), .b(dm_int_st1_28[19]), .cin(dm_int_st1_28[20]), .s(dm_int_st2_28[15]), .cout(dm_int_st2_29[6]));
	full_adder FA58(.a(dm_int_st1_28[21]), .b(dm_int_st1_28[22]), .cin(dm_int_st1_28[23]), .s(dm_int_st2_28[16]), .cout(dm_int_st2_29[7]));
	full_adder FA59(.a(dm_int_st1_28[24]), .b(dm_int_st1_28[25]), .cin(dm_int_st1_28[26]), .s(dm_int_st2_28[17]), .cout(dm_int_st2_29[8]));
	assign dm_int_st2_28[18] = dm_int_st1_28[27];
	// Bit 29
	full_adder FA60(.a(dm_int_st1_29[0]), .b(dm_int_st1_29[1]), .cin(dm_int_st1_29[2]), .s(dm_int_st2_29[9]), .cout(dm_int_st2_30[0]));
	full_adder FA61(.a(dm_int_st1_29[3]), .b(dm_int_st1_29[4]), .cin(dm_int_st1_29[5]), .s(dm_int_st2_29[10]), .cout(dm_int_st2_30[1]));
	full_adder FA62(.a(dm_int_st1_29[6]), .b(dm_int_st1_29[7]), .cin(dm_int_st1_29[8]), .s(dm_int_st2_29[11]), .cout(dm_int_st2_30[2]));
	full_adder FA63(.a(dm_int_st1_29[9]), .b(dm_int_st1_29[10]), .cin(dm_int_st1_29[11]), .s(dm_int_st2_29[12]), .cout(dm_int_st2_30[3]));
	full_adder FA64(.a(dm_int_st1_29[12]), .b(dm_int_st1_29[13]), .cin(dm_int_st1_29[14]), .s(dm_int_st2_29[13]), .cout(dm_int_st2_30[4]));
	full_adder FA65(.a(dm_int_st1_29[15]), .b(dm_int_st1_29[16]), .cin(dm_int_st1_29[17]), .s(dm_int_st2_29[14]), .cout(dm_int_st2_30[5]));
	full_adder FA66(.a(dm_int_st1_29[18]), .b(dm_int_st1_29[19]), .cin(dm_int_st1_29[20]), .s(dm_int_st2_29[15]), .cout(dm_int_st2_30[6]));
	full_adder FA67(.a(dm_int_st1_29[21]), .b(dm_int_st1_29[22]), .cin(dm_int_st1_29[23]), .s(dm_int_st2_29[16]), .cout(dm_int_st2_30[7]));
	full_adder FA68(.a(dm_int_st1_29[24]), .b(dm_int_st1_29[25]), .cin(dm_int_st1_29[26]), .s(dm_int_st2_29[17]), .cout(dm_int_st2_30[8]));
	assign dm_int_st2_29[18] = dm_int_st1_29[27];
	// Bit 30
	full_adder FA69(.a(dm_int_st1_30[0]), .b(dm_int_st1_30[1]), .cin(dm_int_st1_30[2]), .s(dm_int_st2_30[9]), .cout(dm_int_st2_31[0]));
	full_adder FA70(.a(dm_int_st1_30[3]), .b(dm_int_st1_30[4]), .cin(dm_int_st1_30[5]), .s(dm_int_st2_30[10]), .cout(dm_int_st2_31[1]));
	full_adder FA71(.a(dm_int_st1_30[6]), .b(dm_int_st1_30[7]), .cin(dm_int_st1_30[8]), .s(dm_int_st2_30[11]), .cout(dm_int_st2_31[2]));
	full_adder FA72(.a(dm_int_st1_30[9]), .b(dm_int_st1_30[10]), .cin(dm_int_st1_30[11]), .s(dm_int_st2_30[12]), .cout(dm_int_st2_31[3]));
	full_adder FA73(.a(dm_int_st1_30[12]), .b(dm_int_st1_30[13]), .cin(dm_int_st1_30[14]), .s(dm_int_st2_30[13]), .cout(dm_int_st2_31[4]));
	full_adder FA74(.a(dm_int_st1_30[15]), .b(dm_int_st1_30[16]), .cin(dm_int_st1_30[17]), .s(dm_int_st2_30[14]), .cout(dm_int_st2_31[5]));
	full_adder FA75(.a(dm_int_st1_30[18]), .b(dm_int_st1_30[19]), .cin(dm_int_st1_30[20]), .s(dm_int_st2_30[15]), .cout(dm_int_st2_31[6]));
	full_adder FA76(.a(dm_int_st1_30[21]), .b(dm_int_st1_30[22]), .cin(dm_int_st1_30[23]), .s(dm_int_st2_30[16]), .cout(dm_int_st2_31[7]));
	full_adder FA77(.a(dm_int_st1_30[24]), .b(dm_int_st1_30[25]), .cin(dm_int_st1_30[26]), .s(dm_int_st2_30[17]), .cout(dm_int_st2_31[8]));
	assign dm_int_st2_30[18] = dm_int_st1_30[27];
	// Bit 31
	full_adder FA78(.a(dm_int_st1_31[0]), .b(dm_int_st1_31[1]), .cin(dm_int_st1_31[2]), .s(dm_int_st2_31[9]), .cout(dm_int_st2_32[0]));
	full_adder FA79(.a(dm_int_st1_31[3]), .b(dm_int_st1_31[4]), .cin(dm_int_st1_31[5]), .s(dm_int_st2_31[10]), .cout(dm_int_st2_32[1]));
	full_adder FA80(.a(dm_int_st1_31[6]), .b(dm_int_st1_31[7]), .cin(dm_int_st1_31[8]), .s(dm_int_st2_31[11]), .cout(dm_int_st2_32[2]));
	full_adder FA81(.a(dm_int_st1_31[9]), .b(dm_int_st1_31[10]), .cin(dm_int_st1_31[11]), .s(dm_int_st2_31[12]), .cout(dm_int_st2_32[3]));
	full_adder FA82(.a(dm_int_st1_31[12]), .b(dm_int_st1_31[13]), .cin(dm_int_st1_31[14]), .s(dm_int_st2_31[13]), .cout(dm_int_st2_32[4]));
	full_adder FA83(.a(dm_int_st1_31[15]), .b(dm_int_st1_31[16]), .cin(dm_int_st1_31[17]), .s(dm_int_st2_31[14]), .cout(dm_int_st2_32[5]));
	full_adder FA84(.a(dm_int_st1_31[18]), .b(dm_int_st1_31[19]), .cin(dm_int_st1_31[20]), .s(dm_int_st2_31[15]), .cout(dm_int_st2_32[6]));
	full_adder FA85(.a(dm_int_st1_31[21]), .b(dm_int_st1_31[22]), .cin(dm_int_st1_31[23]), .s(dm_int_st2_31[16]), .cout(dm_int_st2_32[7]));
	full_adder FA86(.a(dm_int_st1_31[24]), .b(dm_int_st1_31[25]), .cin(dm_int_st1_31[26]), .s(dm_int_st2_31[17]), .cout(dm_int_st2_32[8]));
	assign dm_int_st2_31[18] = dm_int_st1_31[27];
	// Bit 32
	full_adder FA87(.a(dm_int_st1_32[0]), .b(dm_int_st1_32[1]), .cin(dm_int_st1_32[2]), .s(dm_int_st2_32[9]), .cout(dm_int_st2_33[0]));
	full_adder FA88(.a(dm_int_st1_32[3]), .b(dm_int_st1_32[4]), .cin(dm_int_st1_32[5]), .s(dm_int_st2_32[10]), .cout(dm_int_st2_33[1]));
	full_adder FA89(.a(dm_int_st1_32[6]), .b(dm_int_st1_32[7]), .cin(dm_int_st1_32[8]), .s(dm_int_st2_32[11]), .cout(dm_int_st2_33[2]));
	full_adder FA90(.a(dm_int_st1_32[9]), .b(dm_int_st1_32[10]), .cin(dm_int_st1_32[11]), .s(dm_int_st2_32[12]), .cout(dm_int_st2_33[3]));
	full_adder FA91(.a(dm_int_st1_32[12]), .b(dm_int_st1_32[13]), .cin(dm_int_st1_32[14]), .s(dm_int_st2_32[13]), .cout(dm_int_st2_33[4]));
	full_adder FA92(.a(dm_int_st1_32[15]), .b(dm_int_st1_32[16]), .cin(dm_int_st1_32[17]), .s(dm_int_st2_32[14]), .cout(dm_int_st2_33[5]));
	full_adder FA93(.a(dm_int_st1_32[18]), .b(dm_int_st1_32[19]), .cin(dm_int_st1_32[20]), .s(dm_int_st2_32[15]), .cout(dm_int_st2_33[6]));
	full_adder FA94(.a(dm_int_st1_32[21]), .b(dm_int_st1_32[22]), .cin(dm_int_st1_32[23]), .s(dm_int_st2_32[16]), .cout(dm_int_st2_33[7]));
	full_adder FA95(.a(dm_int_st1_32[24]), .b(dm_int_st1_32[25]), .cin(dm_int_st1_32[26]), .s(dm_int_st2_32[17]), .cout(dm_int_st2_33[8]));
	assign dm_int_st2_32[18] = dm_int_st1_32[27];
	// Bit 33
	full_adder FA96(.a(dm_int_st1_33[0]), .b(dm_int_st1_33[1]), .cin(dm_int_st1_33[2]), .s(dm_int_st2_33[9]), .cout(dm_int_st2_34[0]));
	full_adder FA97(.a(dm_int_st1_33[3]), .b(dm_int_st1_33[4]), .cin(dm_int_st1_33[5]), .s(dm_int_st2_33[10]), .cout(dm_int_st2_34[1]));
	full_adder FA98(.a(dm_int_st1_33[6]), .b(dm_int_st1_33[7]), .cin(dm_int_st1_33[8]), .s(dm_int_st2_33[11]), .cout(dm_int_st2_34[2]));
	full_adder FA99(.a(dm_int_st1_33[9]), .b(dm_int_st1_33[10]), .cin(dm_int_st1_33[11]), .s(dm_int_st2_33[12]), .cout(dm_int_st2_34[3]));
	full_adder FA100(.a(dm_int_st1_33[12]), .b(dm_int_st1_33[13]), .cin(dm_int_st1_33[14]), .s(dm_int_st2_33[13]), .cout(dm_int_st2_34[4]));
	full_adder FA101(.a(dm_int_st1_33[15]), .b(dm_int_st1_33[16]), .cin(dm_int_st1_33[17]), .s(dm_int_st2_33[14]), .cout(dm_int_st2_34[5]));
	full_adder FA102(.a(dm_int_st1_33[18]), .b(dm_int_st1_33[19]), .cin(dm_int_st1_33[20]), .s(dm_int_st2_33[15]), .cout(dm_int_st2_34[6]));
	full_adder FA103(.a(dm_int_st1_33[21]), .b(dm_int_st1_33[22]), .cin(dm_int_st1_33[23]), .s(dm_int_st2_33[16]), .cout(dm_int_st2_34[7]));
	full_adder FA104(.a(dm_int_st1_33[24]), .b(dm_int_st1_33[25]), .cin(dm_int_st1_33[26]), .s(dm_int_st2_33[17]), .cout(dm_int_st2_34[8]));
	assign dm_int_st2_33[18] = dm_int_st1_33[27];
	// Bit 34
	full_adder FA105(.a(dm_int_st1_34[0]), .b(dm_int_st1_34[1]), .cin(dm_int_st1_34[2]), .s(dm_int_st2_34[9]), .cout(dm_int_st2_35[0]));
	full_adder FA106(.a(dm_int_st1_34[3]), .b(dm_int_st1_34[4]), .cin(dm_int_st1_34[5]), .s(dm_int_st2_34[10]), .cout(dm_int_st2_35[1]));
	full_adder FA107(.a(dm_int_st1_34[6]), .b(dm_int_st1_34[7]), .cin(dm_int_st1_34[8]), .s(dm_int_st2_34[11]), .cout(dm_int_st2_35[2]));
	full_adder FA108(.a(dm_int_st1_34[9]), .b(dm_int_st1_34[10]), .cin(dm_int_st1_34[11]), .s(dm_int_st2_34[12]), .cout(dm_int_st2_35[3]));
	full_adder FA109(.a(dm_int_st1_34[12]), .b(dm_int_st1_34[13]), .cin(dm_int_st1_34[14]), .s(dm_int_st2_34[13]), .cout(dm_int_st2_35[4]));
	full_adder FA110(.a(dm_int_st1_34[15]), .b(dm_int_st1_34[16]), .cin(dm_int_st1_34[17]), .s(dm_int_st2_34[14]), .cout(dm_int_st2_35[5]));
	full_adder FA111(.a(dm_int_st1_34[18]), .b(dm_int_st1_34[19]), .cin(dm_int_st1_34[20]), .s(dm_int_st2_34[15]), .cout(dm_int_st2_35[6]));
	full_adder FA112(.a(dm_int_st1_34[21]), .b(dm_int_st1_34[22]), .cin(dm_int_st1_34[23]), .s(dm_int_st2_34[16]), .cout(dm_int_st2_35[7]));
	full_adder FA113(.a(dm_int_st1_34[24]), .b(dm_int_st1_34[25]), .cin(dm_int_st1_34[26]), .s(dm_int_st2_34[17]), .cout(dm_int_st2_35[8]));
	assign dm_int_st2_34[18] = dm_int_st1_34[27];
	// Bit 35
	full_adder FA114(.a(dm_int_st1_35[0]), .b(dm_int_st1_35[1]), .cin(dm_int_st1_35[2]), .s(dm_int_st2_35[9]), .cout(dm_int_st2_36[0]));
	full_adder FA115(.a(dm_int_st1_35[3]), .b(dm_int_st1_35[4]), .cin(dm_int_st1_35[5]), .s(dm_int_st2_35[10]), .cout(dm_int_st2_36[1]));
	full_adder FA116(.a(dm_int_st1_35[6]), .b(dm_int_st1_35[7]), .cin(dm_int_st1_35[8]), .s(dm_int_st2_35[11]), .cout(dm_int_st2_36[2]));
	full_adder FA117(.a(dm_int_st1_35[9]), .b(dm_int_st1_35[10]), .cin(dm_int_st1_35[11]), .s(dm_int_st2_35[12]), .cout(dm_int_st2_36[3]));
	full_adder FA118(.a(dm_int_st1_35[12]), .b(dm_int_st1_35[13]), .cin(dm_int_st1_35[14]), .s(dm_int_st2_35[13]), .cout(dm_int_st2_36[4]));
	full_adder FA119(.a(dm_int_st1_35[15]), .b(dm_int_st1_35[16]), .cin(dm_int_st1_35[17]), .s(dm_int_st2_35[14]), .cout(dm_int_st2_36[5]));
	full_adder FA120(.a(dm_int_st1_35[18]), .b(dm_int_st1_35[19]), .cin(dm_int_st1_35[20]), .s(dm_int_st2_35[15]), .cout(dm_int_st2_36[6]));
	full_adder FA121(.a(dm_int_st1_35[21]), .b(dm_int_st1_35[22]), .cin(dm_int_st1_35[23]), .s(dm_int_st2_35[16]), .cout(dm_int_st2_36[7]));
	full_adder FA122(.a(dm_int_st1_35[24]), .b(dm_int_st1_35[25]), .cin(dm_int_st1_35[26]), .s(dm_int_st2_35[17]), .cout(dm_int_st2_36[8]));
	assign dm_int_st2_35[18] = dm_int_st1_35[27];
	// Bit 36
	full_adder FA123(.a(dm_int_st1_36[0]), .b(dm_int_st1_36[1]), .cin(dm_int_st1_36[2]), .s(dm_int_st2_36[9]), .cout(dm_int_st2_37[0]));
	full_adder FA124(.a(dm_int_st1_36[3]), .b(dm_int_st1_36[4]), .cin(dm_int_st1_36[5]), .s(dm_int_st2_36[10]), .cout(dm_int_st2_37[1]));
	full_adder FA125(.a(dm_int_st1_36[6]), .b(dm_int_st1_36[7]), .cin(dm_int_st1_36[8]), .s(dm_int_st2_36[11]), .cout(dm_int_st2_37[2]));
	full_adder FA126(.a(dm_int_st1_36[9]), .b(dm_int_st1_36[10]), .cin(dm_int_st1_36[11]), .s(dm_int_st2_36[12]), .cout(dm_int_st2_37[3]));
	full_adder FA127(.a(dm_int_st1_36[12]), .b(dm_int_st1_36[13]), .cin(dm_int_st1_36[14]), .s(dm_int_st2_36[13]), .cout(dm_int_st2_37[4]));
	full_adder FA128(.a(dm_int_st1_36[15]), .b(dm_int_st1_36[16]), .cin(dm_int_st1_36[17]), .s(dm_int_st2_36[14]), .cout(dm_int_st2_37[5]));
	full_adder FA129(.a(dm_int_st1_36[18]), .b(dm_int_st1_36[19]), .cin(dm_int_st1_36[20]), .s(dm_int_st2_36[15]), .cout(dm_int_st2_37[6]));
	full_adder FA130(.a(dm_int_st1_36[21]), .b(dm_int_st1_36[22]), .cin(dm_int_st1_36[23]), .s(dm_int_st2_36[16]), .cout(dm_int_st2_37[7]));
	full_adder FA131(.a(dm_int_st1_36[24]), .b(dm_int_st1_36[25]), .cin(dm_int_st1_36[26]), .s(dm_int_st2_36[17]), .cout(dm_int_st2_37[8]));
	assign dm_int_st2_36[18] = dm_int_st1_36[27];
	// Bit 37
	full_adder FA132(.a(dm_int_st1_37[0]), .b(dm_int_st1_37[1]), .cin(dm_int_st1_37[2]), .s(dm_int_st2_37[9]), .cout(dm_int_st2_38[0]));
	full_adder FA133(.a(dm_int_st1_37[3]), .b(dm_int_st1_37[4]), .cin(dm_int_st1_37[5]), .s(dm_int_st2_37[10]), .cout(dm_int_st2_38[1]));
	full_adder FA134(.a(dm_int_st1_37[6]), .b(dm_int_st1_37[7]), .cin(dm_int_st1_37[8]), .s(dm_int_st2_37[11]), .cout(dm_int_st2_38[2]));
	full_adder FA135(.a(dm_int_st1_37[9]), .b(dm_int_st1_37[10]), .cin(dm_int_st1_37[11]), .s(dm_int_st2_37[12]), .cout(dm_int_st2_38[3]));
	full_adder FA136(.a(dm_int_st1_37[12]), .b(dm_int_st1_37[13]), .cin(dm_int_st1_37[14]), .s(dm_int_st2_37[13]), .cout(dm_int_st2_38[4]));
	full_adder FA137(.a(dm_int_st1_37[15]), .b(dm_int_st1_37[16]), .cin(dm_int_st1_37[17]), .s(dm_int_st2_37[14]), .cout(dm_int_st2_38[5]));
	full_adder FA138(.a(dm_int_st1_37[18]), .b(dm_int_st1_37[19]), .cin(dm_int_st1_37[20]), .s(dm_int_st2_37[15]), .cout(dm_int_st2_38[6]));
	full_adder FA139(.a(dm_int_st1_37[21]), .b(dm_int_st1_37[22]), .cin(dm_int_st1_37[23]), .s(dm_int_st2_37[16]), .cout(dm_int_st2_38[7]));
	assign dm_int_st2_37[17] = dm_int_st1_37[24];
	assign dm_int_st2_37[18] = dm_int_st1_37[25];
	// Bit 38
	full_adder FA140(.a(dm_int_st1_38[0]), .b(dm_int_st1_38[1]), .cin(dm_int_st1_38[2]), .s(dm_int_st2_38[8]), .cout(dm_int_st2_39[0]));
	full_adder FA141(.a(dm_int_st1_38[3]), .b(dm_int_st1_38[4]), .cin(dm_int_st1_38[5]), .s(dm_int_st2_38[9]), .cout(dm_int_st2_39[1]));
	full_adder FA142(.a(dm_int_st1_38[6]), .b(dm_int_st1_38[7]), .cin(dm_int_st1_38[8]), .s(dm_int_st2_38[10]), .cout(dm_int_st2_39[2]));
	full_adder FA143(.a(dm_int_st1_38[9]), .b(dm_int_st1_38[10]), .cin(dm_int_st1_38[11]), .s(dm_int_st2_38[11]), .cout(dm_int_st2_39[3]));
	full_adder FA144(.a(dm_int_st1_38[12]), .b(dm_int_st1_38[13]), .cin(dm_int_st1_38[14]), .s(dm_int_st2_38[12]), .cout(dm_int_st2_39[4]));
	full_adder FA145(.a(dm_int_st1_38[15]), .b(dm_int_st1_38[16]), .cin(dm_int_st1_38[17]), .s(dm_int_st2_38[13]), .cout(dm_int_st2_39[5]));
	full_adder FA146(.a(dm_int_st1_38[18]), .b(dm_int_st1_38[19]), .cin(dm_int_st1_38[20]), .s(dm_int_st2_38[14]), .cout(dm_int_st2_39[6]));
	assign dm_int_st2_38[15] = dm_int_st1_38[21];
	assign dm_int_st2_38[16] = dm_int_st1_38[22];
	assign dm_int_st2_38[17] = dm_int_st1_38[23];
	assign dm_int_st2_38[18] = dm_int_st1_38[24];
	// Bit 39
	full_adder FA147(.a(dm_int_st1_39[0]), .b(dm_int_st1_39[1]), .cin(dm_int_st1_39[2]), .s(dm_int_st2_39[7]), .cout(dm_int_st2_40[0]));
	full_adder FA148(.a(dm_int_st1_39[3]), .b(dm_int_st1_39[4]), .cin(dm_int_st1_39[5]), .s(dm_int_st2_39[8]), .cout(dm_int_st2_40[1]));
	full_adder FA149(.a(dm_int_st1_39[6]), .b(dm_int_st1_39[7]), .cin(dm_int_st1_39[8]), .s(dm_int_st2_39[9]), .cout(dm_int_st2_40[2]));
	full_adder FA150(.a(dm_int_st1_39[9]), .b(dm_int_st1_39[10]), .cin(dm_int_st1_39[11]), .s(dm_int_st2_39[10]), .cout(dm_int_st2_40[3]));
	full_adder FA151(.a(dm_int_st1_39[12]), .b(dm_int_st1_39[13]), .cin(dm_int_st1_39[14]), .s(dm_int_st2_39[11]), .cout(dm_int_st2_40[4]));
	full_adder FA152(.a(dm_int_st1_39[15]), .b(dm_int_st1_39[16]), .cin(dm_int_st1_39[17]), .s(dm_int_st2_39[12]), .cout(dm_int_st2_40[5]));
	assign dm_int_st2_39[13] = dm_int_st1_39[18];
	assign dm_int_st2_39[14] = dm_int_st1_39[19];
	assign dm_int_st2_39[15] = dm_int_st1_39[20];
	assign dm_int_st2_39[16] = dm_int_st1_39[21];
	assign dm_int_st2_39[17] = dm_int_st1_39[22];
	assign dm_int_st2_39[18] = dm_int_st1_39[23];
	// Bit 40
	full_adder FA153(.a(dm_int_st1_40[0]), .b(dm_int_st1_40[1]), .cin(dm_int_st1_40[2]), .s(dm_int_st2_40[6]), .cout(dm_int_st2_41[0]));
	full_adder FA154(.a(dm_int_st1_40[3]), .b(dm_int_st1_40[4]), .cin(dm_int_st1_40[5]), .s(dm_int_st2_40[7]), .cout(dm_int_st2_41[1]));
	full_adder FA155(.a(dm_int_st1_40[6]), .b(dm_int_st1_40[7]), .cin(dm_int_st1_40[8]), .s(dm_int_st2_40[8]), .cout(dm_int_st2_41[2]));
	full_adder FA156(.a(dm_int_st1_40[9]), .b(dm_int_st1_40[10]), .cin(dm_int_st1_40[11]), .s(dm_int_st2_40[9]), .cout(dm_int_st2_41[3]));
	full_adder FA157(.a(dm_int_st1_40[12]), .b(dm_int_st1_40[13]), .cin(dm_int_st1_40[14]), .s(dm_int_st2_40[10]), .cout(dm_int_st2_41[4]));
	assign dm_int_st2_40[11] = dm_int_st1_40[15];
	assign dm_int_st2_40[12] = dm_int_st1_40[16];
	assign dm_int_st2_40[13] = dm_int_st1_40[17];
	assign dm_int_st2_40[14] = dm_int_st1_40[18];
	assign dm_int_st2_40[15] = dm_int_st1_40[19];
	assign dm_int_st2_40[16] = dm_int_st1_40[20];
	assign dm_int_st2_40[17] = dm_int_st1_40[21];
	assign dm_int_st2_40[18] = dm_int_st1_40[22];
	// Bit 41
	full_adder FA158(.a(dm_int_st1_41[0]), .b(dm_int_st1_41[1]), .cin(dm_int_st1_41[2]), .s(dm_int_st2_41[5]), .cout(dm_int_st2_42[0]));
	full_adder FA159(.a(dm_int_st1_41[3]), .b(dm_int_st1_41[4]), .cin(dm_int_st1_41[5]), .s(dm_int_st2_41[6]), .cout(dm_int_st2_42[1]));
	full_adder FA160(.a(dm_int_st1_41[6]), .b(dm_int_st1_41[7]), .cin(dm_int_st1_41[8]), .s(dm_int_st2_41[7]), .cout(dm_int_st2_42[2]));
	full_adder FA161(.a(dm_int_st1_41[9]), .b(dm_int_st1_41[10]), .cin(dm_int_st1_41[11]), .s(dm_int_st2_41[8]), .cout(dm_int_st2_42[3]));
	assign dm_int_st2_41[9] = dm_int_st1_41[12];
	assign dm_int_st2_41[10] = dm_int_st1_41[13];
	assign dm_int_st2_41[11] = dm_int_st1_41[14];
	assign dm_int_st2_41[12] = dm_int_st1_41[15];
	assign dm_int_st2_41[13] = dm_int_st1_41[16];
	assign dm_int_st2_41[14] = dm_int_st1_41[17];
	assign dm_int_st2_41[15] = dm_int_st1_41[18];
	assign dm_int_st2_41[16] = dm_int_st1_41[19];
	assign dm_int_st2_41[17] = dm_int_st1_41[20];
	assign dm_int_st2_41[18] = dm_int_st1_41[21];
	// Bit 42
	full_adder FA162(.a(dm_int_st1_42[0]), .b(dm_int_st1_42[1]), .cin(dm_int_st1_42[2]), .s(dm_int_st2_42[4]), .cout(dm_int_st2_43[0]));
	full_adder FA163(.a(dm_int_st1_42[3]), .b(dm_int_st1_42[4]), .cin(dm_int_st1_42[5]), .s(dm_int_st2_42[5]), .cout(dm_int_st2_43[1]));
	full_adder FA164(.a(dm_int_st1_42[6]), .b(dm_int_st1_42[7]), .cin(dm_int_st1_42[8]), .s(dm_int_st2_42[6]), .cout(dm_int_st2_43[2]));
	assign dm_int_st2_42[7] = dm_int_st1_42[9];
	assign dm_int_st2_42[8] = dm_int_st1_42[10];
	assign dm_int_st2_42[9] = dm_int_st1_42[11];
	assign dm_int_st2_42[10] = dm_int_st1_42[12];
	assign dm_int_st2_42[11] = dm_int_st1_42[13];
	assign dm_int_st2_42[12] = dm_int_st1_42[14];
	assign dm_int_st2_42[13] = dm_int_st1_42[15];
	assign dm_int_st2_42[14] = dm_int_st1_42[16];
	assign dm_int_st2_42[15] = dm_int_st1_42[17];
	assign dm_int_st2_42[16] = dm_int_st1_42[18];
	assign dm_int_st2_42[17] = dm_int_st1_42[19];
	assign dm_int_st2_42[18] = dm_int_st1_42[20];
	// Bit 43
	full_adder FA165(.a(dm_int_st1_43[0]), .b(dm_int_st1_43[1]), .cin(dm_int_st1_43[2]), .s(dm_int_st2_43[3]), .cout(dm_int_st2_44[0]));
	full_adder FA166(.a(dm_int_st1_43[3]), .b(dm_int_st1_43[4]), .cin(dm_int_st1_43[5]), .s(dm_int_st2_43[4]), .cout(dm_int_st2_44[1]));
	assign dm_int_st2_43[5] = dm_int_st1_43[6];
	assign dm_int_st2_43[6] = dm_int_st1_43[7];
	assign dm_int_st2_43[7] = dm_int_st1_43[8];
	assign dm_int_st2_43[8] = dm_int_st1_43[9];
	assign dm_int_st2_43[9] = dm_int_st1_43[10];
	assign dm_int_st2_43[10] = dm_int_st1_43[11];
	assign dm_int_st2_43[11] = dm_int_st1_43[12];
	assign dm_int_st2_43[12] = dm_int_st1_43[13];
	assign dm_int_st2_43[13] = dm_int_st1_43[14];
	assign dm_int_st2_43[14] = dm_int_st1_43[15];
	assign dm_int_st2_43[15] = dm_int_st1_43[16];
	assign dm_int_st2_43[16] = dm_int_st1_43[17];
	assign dm_int_st2_43[17] = dm_int_st1_43[18];
	assign dm_int_st2_43[18] = dm_int_st1_43[19];
	// Bit 44
	full_adder FA167(.a(dm_int_st1_44[0]), .b(dm_int_st1_44[1]), .cin(dm_int_st1_44[2]), .s(dm_int_st2_44[2]), .cout(dm_int_st2_45[0]));
	assign dm_int_st2_44[3] = dm_int_st1_44[3];
	assign dm_int_st2_44[4] = dm_int_st1_44[4];
	assign dm_int_st2_44[5] = dm_int_st1_44[5];
	assign dm_int_st2_44[6] = dm_int_st1_44[6];
	assign dm_int_st2_44[7] = dm_int_st1_44[7];
	assign dm_int_st2_44[8] = dm_int_st1_44[8];
	assign dm_int_st2_44[9] = dm_int_st1_44[9];
	assign dm_int_st2_44[10] = dm_int_st1_44[10];
	assign dm_int_st2_44[11] = dm_int_st1_44[11];
	assign dm_int_st2_44[12] = dm_int_st1_44[12];
	assign dm_int_st2_44[13] = dm_int_st1_44[13];
	assign dm_int_st2_44[14] = dm_int_st1_44[14];
	assign dm_int_st2_44[15] = dm_int_st1_44[15];
	assign dm_int_st2_44[16] = dm_int_st1_44[16];
	assign dm_int_st2_44[17] = dm_int_st1_44[17];
	assign dm_int_st2_44[18] = dm_int_st1_44[18];
	// Bit 45
	assign dm_int_st2_45[1] = dm_int_st1_45[0];
	assign dm_int_st2_45[2] = dm_int_st1_45[1];
	assign dm_int_st2_45[3] = dm_int_st1_45[2];
	assign dm_int_st2_45[4] = dm_int_st1_45[3];
	assign dm_int_st2_45[5] = dm_int_st1_45[4];
	assign dm_int_st2_45[6] = dm_int_st1_45[5];
	assign dm_int_st2_45[7] = dm_int_st1_45[6];
	assign dm_int_st2_45[8] = dm_int_st1_45[7];
	assign dm_int_st2_45[9] = dm_int_st1_45[8];
	assign dm_int_st2_45[10] = dm_int_st1_45[9];
	assign dm_int_st2_45[11] = dm_int_st1_45[10];
	assign dm_int_st2_45[12] = dm_int_st1_45[11];
	assign dm_int_st2_45[13] = dm_int_st1_45[12];
	assign dm_int_st2_45[14] = dm_int_st1_45[13];
	assign dm_int_st2_45[15] = dm_int_st1_45[14];
	assign dm_int_st2_45[16] = dm_int_st1_45[15];
	assign dm_int_st2_45[17] = dm_int_st1_45[16];
	assign dm_int_st2_45[18] = dm_int_st1_45[17];
	// Bit 46
	assign dm_int_st2_46[0] = dm_int_st1_46[0];
	assign dm_int_st2_46[1] = dm_int_st1_46[1];
	assign dm_int_st2_46[2] = dm_int_st1_46[2];
	assign dm_int_st2_46[3] = dm_int_st1_46[3];
	assign dm_int_st2_46[4] = dm_int_st1_46[4];
	assign dm_int_st2_46[5] = dm_int_st1_46[5];
	assign dm_int_st2_46[6] = dm_int_st1_46[6];
	assign dm_int_st2_46[7] = dm_int_st1_46[7];
	assign dm_int_st2_46[8] = dm_int_st1_46[8];
	assign dm_int_st2_46[9] = dm_int_st1_46[9];
	assign dm_int_st2_46[10] = dm_int_st1_46[10];
	assign dm_int_st2_46[11] = dm_int_st1_46[11];
	assign dm_int_st2_46[12] = dm_int_st1_46[12];
	assign dm_int_st2_46[13] = dm_int_st1_46[13];
	assign dm_int_st2_46[14] = dm_int_st1_46[14];
	assign dm_int_st2_46[15] = dm_int_st1_46[15];
	assign dm_int_st2_46[16] = dm_int_st1_46[16];
	// Bit 47
	assign dm_int_st2_47[0] = dm_int_st1_47[0];
	assign dm_int_st2_47[1] = dm_int_st1_47[1];
	assign dm_int_st2_47[2] = dm_int_st1_47[2];
	assign dm_int_st2_47[3] = dm_int_st1_47[3];
	assign dm_int_st2_47[4] = dm_int_st1_47[4];
	assign dm_int_st2_47[5] = dm_int_st1_47[5];
	assign dm_int_st2_47[6] = dm_int_st1_47[6];
	assign dm_int_st2_47[7] = dm_int_st1_47[7];
	assign dm_int_st2_47[8] = dm_int_st1_47[8];
	assign dm_int_st2_47[9] = dm_int_st1_47[9];
	assign dm_int_st2_47[10] = dm_int_st1_47[10];
	assign dm_int_st2_47[11] = dm_int_st1_47[11];
	assign dm_int_st2_47[12] = dm_int_st1_47[12];
	assign dm_int_st2_47[13] = dm_int_st1_47[13];
	assign dm_int_st2_47[14] = dm_int_st1_47[14];
	assign dm_int_st2_47[15] = dm_int_st1_47[15];
	// Bit 48
	assign dm_int_st2_48[0] = dm_int_st1_48[0];
	assign dm_int_st2_48[1] = dm_int_st1_48[1];
	assign dm_int_st2_48[2] = dm_int_st1_48[2];
	assign dm_int_st2_48[3] = dm_int_st1_48[3];
	assign dm_int_st2_48[4] = dm_int_st1_48[4];
	assign dm_int_st2_48[5] = dm_int_st1_48[5];
	assign dm_int_st2_48[6] = dm_int_st1_48[6];
	assign dm_int_st2_48[7] = dm_int_st1_48[7];
	assign dm_int_st2_48[8] = dm_int_st1_48[8];
	assign dm_int_st2_48[9] = dm_int_st1_48[9];
	assign dm_int_st2_48[10] = dm_int_st1_48[10];
	assign dm_int_st2_48[11] = dm_int_st1_48[11];
	assign dm_int_st2_48[12] = dm_int_st1_48[12];
	assign dm_int_st2_48[13] = dm_int_st1_48[13];
	assign dm_int_st2_48[14] = dm_int_st1_48[14];
	// Bit 49
	assign dm_int_st2_49[0] = dm_int_st1_49[0];
	assign dm_int_st2_49[1] = dm_int_st1_49[1];
	assign dm_int_st2_49[2] = dm_int_st1_49[2];
	assign dm_int_st2_49[3] = dm_int_st1_49[3];
	assign dm_int_st2_49[4] = dm_int_st1_49[4];
	assign dm_int_st2_49[5] = dm_int_st1_49[5];
	assign dm_int_st2_49[6] = dm_int_st1_49[6];
	assign dm_int_st2_49[7] = dm_int_st1_49[7];
	assign dm_int_st2_49[8] = dm_int_st1_49[8];
	assign dm_int_st2_49[9] = dm_int_st1_49[9];
	assign dm_int_st2_49[10] = dm_int_st1_49[10];
	assign dm_int_st2_49[11] = dm_int_st1_49[11];
	assign dm_int_st2_49[12] = dm_int_st1_49[12];
	assign dm_int_st2_49[13] = dm_int_st1_49[13];
	// Bit 50
	assign dm_int_st2_50[0] = dm_int_st1_50[0];
	assign dm_int_st2_50[1] = dm_int_st1_50[1];
	assign dm_int_st2_50[2] = dm_int_st1_50[2];
	assign dm_int_st2_50[3] = dm_int_st1_50[3];
	assign dm_int_st2_50[4] = dm_int_st1_50[4];
	assign dm_int_st2_50[5] = dm_int_st1_50[5];
	assign dm_int_st2_50[6] = dm_int_st1_50[6];
	assign dm_int_st2_50[7] = dm_int_st1_50[7];
	assign dm_int_st2_50[8] = dm_int_st1_50[8];
	assign dm_int_st2_50[9] = dm_int_st1_50[9];
	assign dm_int_st2_50[10] = dm_int_st1_50[10];
	assign dm_int_st2_50[11] = dm_int_st1_50[11];
	assign dm_int_st2_50[12] = dm_int_st1_50[12];
	// Bit 51
	assign dm_int_st2_51[0] = dm_int_st1_51[0];
	assign dm_int_st2_51[1] = dm_int_st1_51[1];
	assign dm_int_st2_51[2] = dm_int_st1_51[2];
	assign dm_int_st2_51[3] = dm_int_st1_51[3];
	assign dm_int_st2_51[4] = dm_int_st1_51[4];
	assign dm_int_st2_51[5] = dm_int_st1_51[5];
	assign dm_int_st2_51[6] = dm_int_st1_51[6];
	assign dm_int_st2_51[7] = dm_int_st1_51[7];
	assign dm_int_st2_51[8] = dm_int_st1_51[8];
	assign dm_int_st2_51[9] = dm_int_st1_51[9];
	assign dm_int_st2_51[10] = dm_int_st1_51[10];
	assign dm_int_st2_51[11] = dm_int_st1_51[11];
	// Bit 52
	assign dm_int_st2_52[0] = dm_int_st1_52[0];
	assign dm_int_st2_52[1] = dm_int_st1_52[1];
	assign dm_int_st2_52[2] = dm_int_st1_52[2];
	assign dm_int_st2_52[3] = dm_int_st1_52[3];
	assign dm_int_st2_52[4] = dm_int_st1_52[4];
	assign dm_int_st2_52[5] = dm_int_st1_52[5];
	assign dm_int_st2_52[6] = dm_int_st1_52[6];
	assign dm_int_st2_52[7] = dm_int_st1_52[7];
	assign dm_int_st2_52[8] = dm_int_st1_52[8];
	assign dm_int_st2_52[9] = dm_int_st1_52[9];
	assign dm_int_st2_52[10] = dm_int_st1_52[10];
	// Bit 53
	assign dm_int_st2_53[0] = dm_int_st1_53[0];
	assign dm_int_st2_53[1] = dm_int_st1_53[1];
	assign dm_int_st2_53[2] = dm_int_st1_53[2];
	assign dm_int_st2_53[3] = dm_int_st1_53[3];
	assign dm_int_st2_53[4] = dm_int_st1_53[4];
	assign dm_int_st2_53[5] = dm_int_st1_53[5];
	assign dm_int_st2_53[6] = dm_int_st1_53[6];
	assign dm_int_st2_53[7] = dm_int_st1_53[7];
	assign dm_int_st2_53[8] = dm_int_st1_53[8];
	assign dm_int_st2_53[9] = dm_int_st1_53[9];
	// Bit 54
	assign dm_int_st2_54[0] = dm_int_st1_54[0];
	assign dm_int_st2_54[1] = dm_int_st1_54[1];
	assign dm_int_st2_54[2] = dm_int_st1_54[2];
	assign dm_int_st2_54[3] = dm_int_st1_54[3];
	assign dm_int_st2_54[4] = dm_int_st1_54[4];
	assign dm_int_st2_54[5] = dm_int_st1_54[5];
	assign dm_int_st2_54[6] = dm_int_st1_54[6];
	assign dm_int_st2_54[7] = dm_int_st1_54[7];
	assign dm_int_st2_54[8] = dm_int_st1_54[8];
	// Bit 55
	assign dm_int_st2_55[0] = dm_int_st1_55[0];
	assign dm_int_st2_55[1] = dm_int_st1_55[1];
	assign dm_int_st2_55[2] = dm_int_st1_55[2];
	assign dm_int_st2_55[3] = dm_int_st1_55[3];
	assign dm_int_st2_55[4] = dm_int_st1_55[4];
	assign dm_int_st2_55[5] = dm_int_st1_55[5];
	assign dm_int_st2_55[6] = dm_int_st1_55[6];
	assign dm_int_st2_55[7] = dm_int_st1_55[7];
	// Bit 56
	assign dm_int_st2_56[0] = dm_int_st1_56[0];
	assign dm_int_st2_56[1] = dm_int_st1_56[1];
	assign dm_int_st2_56[2] = dm_int_st1_56[2];
	assign dm_int_st2_56[3] = dm_int_st1_56[3];
	assign dm_int_st2_56[4] = dm_int_st1_56[4];
	assign dm_int_st2_56[5] = dm_int_st1_56[5];
	assign dm_int_st2_56[6] = dm_int_st1_56[6];
	// Bit 57
	assign dm_int_st2_57[0] = dm_int_st1_57[0];
	assign dm_int_st2_57[1] = dm_int_st1_57[1];
	assign dm_int_st2_57[2] = dm_int_st1_57[2];
	assign dm_int_st2_57[3] = dm_int_st1_57[3];
	assign dm_int_st2_57[4] = dm_int_st1_57[4];
	assign dm_int_st2_57[5] = dm_int_st1_57[5];
	// Bit 58
	assign dm_int_st2_58[0] = dm_int_st1_58[0];
	assign dm_int_st2_58[1] = dm_int_st1_58[1];
	assign dm_int_st2_58[2] = dm_int_st1_58[2];
	assign dm_int_st2_58[3] = dm_int_st1_58[3];
	assign dm_int_st2_58[4] = dm_int_st1_58[4];
	// Bit 59
	assign dm_int_st2_59[0] = dm_int_st1_59[0];
	assign dm_int_st2_59[1] = dm_int_st1_59[1];
	assign dm_int_st2_59[2] = dm_int_st1_59[2];
	assign dm_int_st2_59[3] = dm_int_st1_59[3];
	// Bit 60
	assign dm_int_st2_60[0] = dm_int_st1_60[0];
	assign dm_int_st2_60[1] = dm_int_st1_60[1];
	assign dm_int_st2_60[2] = dm_int_st1_60[2];
	// Bit 61
	assign dm_int_st2_61[0] = dm_int_st1_61[0];
	assign dm_int_st2_61[1] = dm_int_st1_61[1];
	// Bit 62
	assign dm_int_st2_62[0] = dm_int_st1_62[0];

	//// Stage 3 ////
	wire [0:0] dm_int_st3_0;
	wire [1:0] dm_int_st3_1;
	wire [2:0] dm_int_st3_2;
	wire [3:0] dm_int_st3_3;
	wire [4:0] dm_int_st3_4;
	wire [5:0] dm_int_st3_5;
	wire [6:0] dm_int_st3_6;
	wire [7:0] dm_int_st3_7;
	wire [8:0] dm_int_st3_8;
	wire [9:0] dm_int_st3_9;
	wire [10:0] dm_int_st3_10;
	wire [11:0] dm_int_st3_11;
	wire [12:0] dm_int_st3_12;
	wire [12:0] dm_int_st3_13;
	wire [12:0] dm_int_st3_14;
	wire [12:0] dm_int_st3_15;
	wire [12:0] dm_int_st3_16;
	wire [12:0] dm_int_st3_17;
	wire [12:0] dm_int_st3_18;
	wire [12:0] dm_int_st3_19;
	wire [12:0] dm_int_st3_20;
	wire [12:0] dm_int_st3_21;
	wire [12:0] dm_int_st3_22;
	wire [12:0] dm_int_st3_23;
	wire [12:0] dm_int_st3_24;
	wire [12:0] dm_int_st3_25;
	wire [12:0] dm_int_st3_26;
	wire [12:0] dm_int_st3_27;
	wire [12:0] dm_int_st3_28;
	wire [12:0] dm_int_st3_29;
	wire [12:0] dm_int_st3_30;
	wire [12:0] dm_int_st3_31;
	wire [12:0] dm_int_st3_32;
	wire [12:0] dm_int_st3_33;
	wire [12:0] dm_int_st3_34;
	wire [12:0] dm_int_st3_35;
	wire [12:0] dm_int_st3_36;
	wire [12:0] dm_int_st3_37;
	wire [12:0] dm_int_st3_38;
	wire [12:0] dm_int_st3_39;
	wire [12:0] dm_int_st3_40;
	wire [12:0] dm_int_st3_41;
	wire [12:0] dm_int_st3_42;
	wire [12:0] dm_int_st3_43;
	wire [12:0] dm_int_st3_44;
	wire [12:0] dm_int_st3_45;
	wire [12:0] dm_int_st3_46;
	wire [12:0] dm_int_st3_47;
	wire [12:0] dm_int_st3_48;
	wire [12:0] dm_int_st3_49;
	wire [12:0] dm_int_st3_50;
	wire [12:0] dm_int_st3_51;
	wire [10:0] dm_int_st3_52;
	wire [9:0] dm_int_st3_53;
	wire [8:0] dm_int_st3_54;
	wire [7:0] dm_int_st3_55;
	wire [6:0] dm_int_st3_56;
	wire [5:0] dm_int_st3_57;
	wire [4:0] dm_int_st3_58;
	wire [3:0] dm_int_st3_59;
	wire [2:0] dm_int_st3_60;
	wire [1:0] dm_int_st3_61;
	wire [0:0] dm_int_st3_62;

	// Bit 0
	assign dm_int_st3_0[0] = dm_int_st2_0[0];
	// Bit 1
	assign dm_int_st3_1[0] = dm_int_st2_1[0];
	assign dm_int_st3_1[1] = dm_int_st2_1[1];
	// Bit 2
	assign dm_int_st3_2[0] = dm_int_st2_2[0];
	assign dm_int_st3_2[1] = dm_int_st2_2[1];
	assign dm_int_st3_2[2] = dm_int_st2_2[2];
	// Bit 3
	assign dm_int_st3_3[0] = dm_int_st2_3[0];
	assign dm_int_st3_3[1] = dm_int_st2_3[1];
	assign dm_int_st3_3[2] = dm_int_st2_3[2];
	assign dm_int_st3_3[3] = dm_int_st2_3[3];
	// Bit 4
	assign dm_int_st3_4[0] = dm_int_st2_4[0];
	assign dm_int_st3_4[1] = dm_int_st2_4[1];
	assign dm_int_st3_4[2] = dm_int_st2_4[2];
	assign dm_int_st3_4[3] = dm_int_st2_4[3];
	assign dm_int_st3_4[4] = dm_int_st2_4[4];
	// Bit 5
	assign dm_int_st3_5[0] = dm_int_st2_5[0];
	assign dm_int_st3_5[1] = dm_int_st2_5[1];
	assign dm_int_st3_5[2] = dm_int_st2_5[2];
	assign dm_int_st3_5[3] = dm_int_st2_5[3];
	assign dm_int_st3_5[4] = dm_int_st2_5[4];
	assign dm_int_st3_5[5] = dm_int_st2_5[5];
	// Bit 6
	assign dm_int_st3_6[0] = dm_int_st2_6[0];
	assign dm_int_st3_6[1] = dm_int_st2_6[1];
	assign dm_int_st3_6[2] = dm_int_st2_6[2];
	assign dm_int_st3_6[3] = dm_int_st2_6[3];
	assign dm_int_st3_6[4] = dm_int_st2_6[4];
	assign dm_int_st3_6[5] = dm_int_st2_6[5];
	assign dm_int_st3_6[6] = dm_int_st2_6[6];
	// Bit 7
	assign dm_int_st3_7[0] = dm_int_st2_7[0];
	assign dm_int_st3_7[1] = dm_int_st2_7[1];
	assign dm_int_st3_7[2] = dm_int_st2_7[2];
	assign dm_int_st3_7[3] = dm_int_st2_7[3];
	assign dm_int_st3_7[4] = dm_int_st2_7[4];
	assign dm_int_st3_7[5] = dm_int_st2_7[5];
	assign dm_int_st3_7[6] = dm_int_st2_7[6];
	assign dm_int_st3_7[7] = dm_int_st2_7[7];
	// Bit 8
	assign dm_int_st3_8[0] = dm_int_st2_8[0];
	assign dm_int_st3_8[1] = dm_int_st2_8[1];
	assign dm_int_st3_8[2] = dm_int_st2_8[2];
	assign dm_int_st3_8[3] = dm_int_st2_8[3];
	assign dm_int_st3_8[4] = dm_int_st2_8[4];
	assign dm_int_st3_8[5] = dm_int_st2_8[5];
	assign dm_int_st3_8[6] = dm_int_st2_8[6];
	assign dm_int_st3_8[7] = dm_int_st2_8[7];
	assign dm_int_st3_8[8] = dm_int_st2_8[8];
	// Bit 9
	assign dm_int_st3_9[0] = dm_int_st2_9[0];
	assign dm_int_st3_9[1] = dm_int_st2_9[1];
	assign dm_int_st3_9[2] = dm_int_st2_9[2];
	assign dm_int_st3_9[3] = dm_int_st2_9[3];
	assign dm_int_st3_9[4] = dm_int_st2_9[4];
	assign dm_int_st3_9[5] = dm_int_st2_9[5];
	assign dm_int_st3_9[6] = dm_int_st2_9[6];
	assign dm_int_st3_9[7] = dm_int_st2_9[7];
	assign dm_int_st3_9[8] = dm_int_st2_9[8];
	assign dm_int_st3_9[9] = dm_int_st2_9[9];
	// Bit 10
	assign dm_int_st3_10[0] = dm_int_st2_10[0];
	assign dm_int_st3_10[1] = dm_int_st2_10[1];
	assign dm_int_st3_10[2] = dm_int_st2_10[2];
	assign dm_int_st3_10[3] = dm_int_st2_10[3];
	assign dm_int_st3_10[4] = dm_int_st2_10[4];
	assign dm_int_st3_10[5] = dm_int_st2_10[5];
	assign dm_int_st3_10[6] = dm_int_st2_10[6];
	assign dm_int_st3_10[7] = dm_int_st2_10[7];
	assign dm_int_st3_10[8] = dm_int_st2_10[8];
	assign dm_int_st3_10[9] = dm_int_st2_10[9];
	assign dm_int_st3_10[10] = dm_int_st2_10[10];
	// Bit 11
	assign dm_int_st3_11[0] = dm_int_st2_11[0];
	assign dm_int_st3_11[1] = dm_int_st2_11[1];
	assign dm_int_st3_11[2] = dm_int_st2_11[2];
	assign dm_int_st3_11[3] = dm_int_st2_11[3];
	assign dm_int_st3_11[4] = dm_int_st2_11[4];
	assign dm_int_st3_11[5] = dm_int_st2_11[5];
	assign dm_int_st3_11[6] = dm_int_st2_11[6];
	assign dm_int_st3_11[7] = dm_int_st2_11[7];
	assign dm_int_st3_11[8] = dm_int_st2_11[8];
	assign dm_int_st3_11[9] = dm_int_st2_11[9];
	assign dm_int_st3_11[10] = dm_int_st2_11[10];
	assign dm_int_st3_11[11] = dm_int_st2_11[11];
	// Bit 12
	assign dm_int_st3_12[0] = dm_int_st2_12[0];
	assign dm_int_st3_12[1] = dm_int_st2_12[1];
	assign dm_int_st3_12[2] = dm_int_st2_12[2];
	assign dm_int_st3_12[3] = dm_int_st2_12[3];
	assign dm_int_st3_12[4] = dm_int_st2_12[4];
	assign dm_int_st3_12[5] = dm_int_st2_12[5];
	assign dm_int_st3_12[6] = dm_int_st2_12[6];
	assign dm_int_st3_12[7] = dm_int_st2_12[7];
	assign dm_int_st3_12[8] = dm_int_st2_12[8];
	assign dm_int_st3_12[9] = dm_int_st2_12[9];
	assign dm_int_st3_12[10] = dm_int_st2_12[10];
	assign dm_int_st3_12[11] = dm_int_st2_12[11];
	assign dm_int_st3_12[12] = dm_int_st2_12[12];
	// Bit 13
	half_adder HA14(.a(dm_int_st2_13[0]), .b(dm_int_st2_13[1]), .s(dm_int_st3_13[0]), .cout(dm_int_st3_14[0]));
	assign dm_int_st3_13[1] = dm_int_st2_13[2];
	assign dm_int_st3_13[2] = dm_int_st2_13[3];
	assign dm_int_st3_13[3] = dm_int_st2_13[4];
	assign dm_int_st3_13[4] = dm_int_st2_13[5];
	assign dm_int_st3_13[5] = dm_int_st2_13[6];
	assign dm_int_st3_13[6] = dm_int_st2_13[7];
	assign dm_int_st3_13[7] = dm_int_st2_13[8];
	assign dm_int_st3_13[8] = dm_int_st2_13[9];
	assign dm_int_st3_13[9] = dm_int_st2_13[10];
	assign dm_int_st3_13[10] = dm_int_st2_13[11];
	assign dm_int_st3_13[11] = dm_int_st2_13[12];
	assign dm_int_st3_13[12] = dm_int_st2_13[13];
	// Bit 14
	full_adder FA168(.a(dm_int_st2_14[0]), .b(dm_int_st2_14[1]), .cin(dm_int_st2_14[2]), .s(dm_int_st3_14[1]), .cout(dm_int_st3_15[0]));
	half_adder HA15(.a(dm_int_st2_14[3]), .b(dm_int_st2_14[4]), .s(dm_int_st3_14[2]), .cout(dm_int_st3_15[1]));
	assign dm_int_st3_14[3] = dm_int_st2_14[5];
	assign dm_int_st3_14[4] = dm_int_st2_14[6];
	assign dm_int_st3_14[5] = dm_int_st2_14[7];
	assign dm_int_st3_14[6] = dm_int_st2_14[8];
	assign dm_int_st3_14[7] = dm_int_st2_14[9];
	assign dm_int_st3_14[8] = dm_int_st2_14[10];
	assign dm_int_st3_14[9] = dm_int_st2_14[11];
	assign dm_int_st3_14[10] = dm_int_st2_14[12];
	assign dm_int_st3_14[11] = dm_int_st2_14[13];
	assign dm_int_st3_14[12] = dm_int_st2_14[14];
	// Bit 15
	full_adder FA169(.a(dm_int_st2_15[0]), .b(dm_int_st2_15[1]), .cin(dm_int_st2_15[2]), .s(dm_int_st3_15[2]), .cout(dm_int_st3_16[0]));
	full_adder FA170(.a(dm_int_st2_15[3]), .b(dm_int_st2_15[4]), .cin(dm_int_st2_15[5]), .s(dm_int_st3_15[3]), .cout(dm_int_st3_16[1]));
	half_adder HA16(.a(dm_int_st2_15[6]), .b(dm_int_st2_15[7]), .s(dm_int_st3_15[4]), .cout(dm_int_st3_16[2]));
	assign dm_int_st3_15[5] = dm_int_st2_15[8];
	assign dm_int_st3_15[6] = dm_int_st2_15[9];
	assign dm_int_st3_15[7] = dm_int_st2_15[10];
	assign dm_int_st3_15[8] = dm_int_st2_15[11];
	assign dm_int_st3_15[9] = dm_int_st2_15[12];
	assign dm_int_st3_15[10] = dm_int_st2_15[13];
	assign dm_int_st3_15[11] = dm_int_st2_15[14];
	assign dm_int_st3_15[12] = dm_int_st2_15[15];
	// Bit 16
	full_adder FA171(.a(dm_int_st2_16[0]), .b(dm_int_st2_16[1]), .cin(dm_int_st2_16[2]), .s(dm_int_st3_16[3]), .cout(dm_int_st3_17[0]));
	full_adder FA172(.a(dm_int_st2_16[3]), .b(dm_int_st2_16[4]), .cin(dm_int_st2_16[5]), .s(dm_int_st3_16[4]), .cout(dm_int_st3_17[1]));
	full_adder FA173(.a(dm_int_st2_16[6]), .b(dm_int_st2_16[7]), .cin(dm_int_st2_16[8]), .s(dm_int_st3_16[5]), .cout(dm_int_st3_17[2]));
	half_adder HA17(.a(dm_int_st2_16[9]), .b(dm_int_st2_16[10]), .s(dm_int_st3_16[6]), .cout(dm_int_st3_17[3]));
	assign dm_int_st3_16[7] = dm_int_st2_16[11];
	assign dm_int_st3_16[8] = dm_int_st2_16[12];
	assign dm_int_st3_16[9] = dm_int_st2_16[13];
	assign dm_int_st3_16[10] = dm_int_st2_16[14];
	assign dm_int_st3_16[11] = dm_int_st2_16[15];
	assign dm_int_st3_16[12] = dm_int_st2_16[16];
	// Bit 17
	full_adder FA174(.a(dm_int_st2_17[0]), .b(dm_int_st2_17[1]), .cin(dm_int_st2_17[2]), .s(dm_int_st3_17[4]), .cout(dm_int_st3_18[0]));
	full_adder FA175(.a(dm_int_st2_17[3]), .b(dm_int_st2_17[4]), .cin(dm_int_st2_17[5]), .s(dm_int_st3_17[5]), .cout(dm_int_st3_18[1]));
	full_adder FA176(.a(dm_int_st2_17[6]), .b(dm_int_st2_17[7]), .cin(dm_int_st2_17[8]), .s(dm_int_st3_17[6]), .cout(dm_int_st3_18[2]));
	full_adder FA177(.a(dm_int_st2_17[9]), .b(dm_int_st2_17[10]), .cin(dm_int_st2_17[11]), .s(dm_int_st3_17[7]), .cout(dm_int_st3_18[3]));
	half_adder HA18(.a(dm_int_st2_17[12]), .b(dm_int_st2_17[13]), .s(dm_int_st3_17[8]), .cout(dm_int_st3_18[4]));
	assign dm_int_st3_17[9] = dm_int_st2_17[14];
	assign dm_int_st3_17[10] = dm_int_st2_17[15];
	assign dm_int_st3_17[11] = dm_int_st2_17[16];
	assign dm_int_st3_17[12] = dm_int_st2_17[17];
	// Bit 18
	full_adder FA178(.a(dm_int_st2_18[0]), .b(dm_int_st2_18[1]), .cin(dm_int_st2_18[2]), .s(dm_int_st3_18[5]), .cout(dm_int_st3_19[0]));
	full_adder FA179(.a(dm_int_st2_18[3]), .b(dm_int_st2_18[4]), .cin(dm_int_st2_18[5]), .s(dm_int_st3_18[6]), .cout(dm_int_st3_19[1]));
	full_adder FA180(.a(dm_int_st2_18[6]), .b(dm_int_st2_18[7]), .cin(dm_int_st2_18[8]), .s(dm_int_st3_18[7]), .cout(dm_int_st3_19[2]));
	full_adder FA181(.a(dm_int_st2_18[9]), .b(dm_int_st2_18[10]), .cin(dm_int_st2_18[11]), .s(dm_int_st3_18[8]), .cout(dm_int_st3_19[3]));
	full_adder FA182(.a(dm_int_st2_18[12]), .b(dm_int_st2_18[13]), .cin(dm_int_st2_18[14]), .s(dm_int_st3_18[9]), .cout(dm_int_st3_19[4]));
	half_adder HA19(.a(dm_int_st2_18[15]), .b(dm_int_st2_18[16]), .s(dm_int_st3_18[10]), .cout(dm_int_st3_19[5]));
	assign dm_int_st3_18[11] = dm_int_st2_18[17];
	assign dm_int_st3_18[12] = dm_int_st2_18[18];
	// Bit 19
	full_adder FA183(.a(dm_int_st2_19[0]), .b(dm_int_st2_19[1]), .cin(dm_int_st2_19[2]), .s(dm_int_st3_19[6]), .cout(dm_int_st3_20[0]));
	full_adder FA184(.a(dm_int_st2_19[3]), .b(dm_int_st2_19[4]), .cin(dm_int_st2_19[5]), .s(dm_int_st3_19[7]), .cout(dm_int_st3_20[1]));
	full_adder FA185(.a(dm_int_st2_19[6]), .b(dm_int_st2_19[7]), .cin(dm_int_st2_19[8]), .s(dm_int_st3_19[8]), .cout(dm_int_st3_20[2]));
	full_adder FA186(.a(dm_int_st2_19[9]), .b(dm_int_st2_19[10]), .cin(dm_int_st2_19[11]), .s(dm_int_st3_19[9]), .cout(dm_int_st3_20[3]));
	full_adder FA187(.a(dm_int_st2_19[12]), .b(dm_int_st2_19[13]), .cin(dm_int_st2_19[14]), .s(dm_int_st3_19[10]), .cout(dm_int_st3_20[4]));
	full_adder FA188(.a(dm_int_st2_19[15]), .b(dm_int_st2_19[16]), .cin(dm_int_st2_19[17]), .s(dm_int_st3_19[11]), .cout(dm_int_st3_20[5]));
	assign dm_int_st3_19[12] = dm_int_st2_19[18];
	// Bit 20
	full_adder FA189(.a(dm_int_st2_20[0]), .b(dm_int_st2_20[1]), .cin(dm_int_st2_20[2]), .s(dm_int_st3_20[6]), .cout(dm_int_st3_21[0]));
	full_adder FA190(.a(dm_int_st2_20[3]), .b(dm_int_st2_20[4]), .cin(dm_int_st2_20[5]), .s(dm_int_st3_20[7]), .cout(dm_int_st3_21[1]));
	full_adder FA191(.a(dm_int_st2_20[6]), .b(dm_int_st2_20[7]), .cin(dm_int_st2_20[8]), .s(dm_int_st3_20[8]), .cout(dm_int_st3_21[2]));
	full_adder FA192(.a(dm_int_st2_20[9]), .b(dm_int_st2_20[10]), .cin(dm_int_st2_20[11]), .s(dm_int_st3_20[9]), .cout(dm_int_st3_21[3]));
	full_adder FA193(.a(dm_int_st2_20[12]), .b(dm_int_st2_20[13]), .cin(dm_int_st2_20[14]), .s(dm_int_st3_20[10]), .cout(dm_int_st3_21[4]));
	full_adder FA194(.a(dm_int_st2_20[15]), .b(dm_int_st2_20[16]), .cin(dm_int_st2_20[17]), .s(dm_int_st3_20[11]), .cout(dm_int_st3_21[5]));
	assign dm_int_st3_20[12] = dm_int_st2_20[18];
	// Bit 21
	full_adder FA195(.a(dm_int_st2_21[0]), .b(dm_int_st2_21[1]), .cin(dm_int_st2_21[2]), .s(dm_int_st3_21[6]), .cout(dm_int_st3_22[0]));
	full_adder FA196(.a(dm_int_st2_21[3]), .b(dm_int_st2_21[4]), .cin(dm_int_st2_21[5]), .s(dm_int_st3_21[7]), .cout(dm_int_st3_22[1]));
	full_adder FA197(.a(dm_int_st2_21[6]), .b(dm_int_st2_21[7]), .cin(dm_int_st2_21[8]), .s(dm_int_st3_21[8]), .cout(dm_int_st3_22[2]));
	full_adder FA198(.a(dm_int_st2_21[9]), .b(dm_int_st2_21[10]), .cin(dm_int_st2_21[11]), .s(dm_int_st3_21[9]), .cout(dm_int_st3_22[3]));
	full_adder FA199(.a(dm_int_st2_21[12]), .b(dm_int_st2_21[13]), .cin(dm_int_st2_21[14]), .s(dm_int_st3_21[10]), .cout(dm_int_st3_22[4]));
	full_adder FA200(.a(dm_int_st2_21[15]), .b(dm_int_st2_21[16]), .cin(dm_int_st2_21[17]), .s(dm_int_st3_21[11]), .cout(dm_int_st3_22[5]));
	assign dm_int_st3_21[12] = dm_int_st2_21[18];
	// Bit 22
	full_adder FA201(.a(dm_int_st2_22[0]), .b(dm_int_st2_22[1]), .cin(dm_int_st2_22[2]), .s(dm_int_st3_22[6]), .cout(dm_int_st3_23[0]));
	full_adder FA202(.a(dm_int_st2_22[3]), .b(dm_int_st2_22[4]), .cin(dm_int_st2_22[5]), .s(dm_int_st3_22[7]), .cout(dm_int_st3_23[1]));
	full_adder FA203(.a(dm_int_st2_22[6]), .b(dm_int_st2_22[7]), .cin(dm_int_st2_22[8]), .s(dm_int_st3_22[8]), .cout(dm_int_st3_23[2]));
	full_adder FA204(.a(dm_int_st2_22[9]), .b(dm_int_st2_22[10]), .cin(dm_int_st2_22[11]), .s(dm_int_st3_22[9]), .cout(dm_int_st3_23[3]));
	full_adder FA205(.a(dm_int_st2_22[12]), .b(dm_int_st2_22[13]), .cin(dm_int_st2_22[14]), .s(dm_int_st3_22[10]), .cout(dm_int_st3_23[4]));
	full_adder FA206(.a(dm_int_st2_22[15]), .b(dm_int_st2_22[16]), .cin(dm_int_st2_22[17]), .s(dm_int_st3_22[11]), .cout(dm_int_st3_23[5]));
	assign dm_int_st3_22[12] = dm_int_st2_22[18];
	// Bit 23
	full_adder FA207(.a(dm_int_st2_23[0]), .b(dm_int_st2_23[1]), .cin(dm_int_st2_23[2]), .s(dm_int_st3_23[6]), .cout(dm_int_st3_24[0]));
	full_adder FA208(.a(dm_int_st2_23[3]), .b(dm_int_st2_23[4]), .cin(dm_int_st2_23[5]), .s(dm_int_st3_23[7]), .cout(dm_int_st3_24[1]));
	full_adder FA209(.a(dm_int_st2_23[6]), .b(dm_int_st2_23[7]), .cin(dm_int_st2_23[8]), .s(dm_int_st3_23[8]), .cout(dm_int_st3_24[2]));
	full_adder FA210(.a(dm_int_st2_23[9]), .b(dm_int_st2_23[10]), .cin(dm_int_st2_23[11]), .s(dm_int_st3_23[9]), .cout(dm_int_st3_24[3]));
	full_adder FA211(.a(dm_int_st2_23[12]), .b(dm_int_st2_23[13]), .cin(dm_int_st2_23[14]), .s(dm_int_st3_23[10]), .cout(dm_int_st3_24[4]));
	full_adder FA212(.a(dm_int_st2_23[15]), .b(dm_int_st2_23[16]), .cin(dm_int_st2_23[17]), .s(dm_int_st3_23[11]), .cout(dm_int_st3_24[5]));
	assign dm_int_st3_23[12] = dm_int_st2_23[18];
	// Bit 24
	full_adder FA213(.a(dm_int_st2_24[0]), .b(dm_int_st2_24[1]), .cin(dm_int_st2_24[2]), .s(dm_int_st3_24[6]), .cout(dm_int_st3_25[0]));
	full_adder FA214(.a(dm_int_st2_24[3]), .b(dm_int_st2_24[4]), .cin(dm_int_st2_24[5]), .s(dm_int_st3_24[7]), .cout(dm_int_st3_25[1]));
	full_adder FA215(.a(dm_int_st2_24[6]), .b(dm_int_st2_24[7]), .cin(dm_int_st2_24[8]), .s(dm_int_st3_24[8]), .cout(dm_int_st3_25[2]));
	full_adder FA216(.a(dm_int_st2_24[9]), .b(dm_int_st2_24[10]), .cin(dm_int_st2_24[11]), .s(dm_int_st3_24[9]), .cout(dm_int_st3_25[3]));
	full_adder FA217(.a(dm_int_st2_24[12]), .b(dm_int_st2_24[13]), .cin(dm_int_st2_24[14]), .s(dm_int_st3_24[10]), .cout(dm_int_st3_25[4]));
	full_adder FA218(.a(dm_int_st2_24[15]), .b(dm_int_st2_24[16]), .cin(dm_int_st2_24[17]), .s(dm_int_st3_24[11]), .cout(dm_int_st3_25[5]));
	assign dm_int_st3_24[12] = dm_int_st2_24[18];
	// Bit 25
	full_adder FA219(.a(dm_int_st2_25[0]), .b(dm_int_st2_25[1]), .cin(dm_int_st2_25[2]), .s(dm_int_st3_25[6]), .cout(dm_int_st3_26[0]));
	full_adder FA220(.a(dm_int_st2_25[3]), .b(dm_int_st2_25[4]), .cin(dm_int_st2_25[5]), .s(dm_int_st3_25[7]), .cout(dm_int_st3_26[1]));
	full_adder FA221(.a(dm_int_st2_25[6]), .b(dm_int_st2_25[7]), .cin(dm_int_st2_25[8]), .s(dm_int_st3_25[8]), .cout(dm_int_st3_26[2]));
	full_adder FA222(.a(dm_int_st2_25[9]), .b(dm_int_st2_25[10]), .cin(dm_int_st2_25[11]), .s(dm_int_st3_25[9]), .cout(dm_int_st3_26[3]));
	full_adder FA223(.a(dm_int_st2_25[12]), .b(dm_int_st2_25[13]), .cin(dm_int_st2_25[14]), .s(dm_int_st3_25[10]), .cout(dm_int_st3_26[4]));
	full_adder FA224(.a(dm_int_st2_25[15]), .b(dm_int_st2_25[16]), .cin(dm_int_st2_25[17]), .s(dm_int_st3_25[11]), .cout(dm_int_st3_26[5]));
	assign dm_int_st3_25[12] = dm_int_st2_25[18];
	// Bit 26
	full_adder FA225(.a(dm_int_st2_26[0]), .b(dm_int_st2_26[1]), .cin(dm_int_st2_26[2]), .s(dm_int_st3_26[6]), .cout(dm_int_st3_27[0]));
	full_adder FA226(.a(dm_int_st2_26[3]), .b(dm_int_st2_26[4]), .cin(dm_int_st2_26[5]), .s(dm_int_st3_26[7]), .cout(dm_int_st3_27[1]));
	full_adder FA227(.a(dm_int_st2_26[6]), .b(dm_int_st2_26[7]), .cin(dm_int_st2_26[8]), .s(dm_int_st3_26[8]), .cout(dm_int_st3_27[2]));
	full_adder FA228(.a(dm_int_st2_26[9]), .b(dm_int_st2_26[10]), .cin(dm_int_st2_26[11]), .s(dm_int_st3_26[9]), .cout(dm_int_st3_27[3]));
	full_adder FA229(.a(dm_int_st2_26[12]), .b(dm_int_st2_26[13]), .cin(dm_int_st2_26[14]), .s(dm_int_st3_26[10]), .cout(dm_int_st3_27[4]));
	full_adder FA230(.a(dm_int_st2_26[15]), .b(dm_int_st2_26[16]), .cin(dm_int_st2_26[17]), .s(dm_int_st3_26[11]), .cout(dm_int_st3_27[5]));
	assign dm_int_st3_26[12] = dm_int_st2_26[18];
	// Bit 27
	full_adder FA231(.a(dm_int_st2_27[0]), .b(dm_int_st2_27[1]), .cin(dm_int_st2_27[2]), .s(dm_int_st3_27[6]), .cout(dm_int_st3_28[0]));
	full_adder FA232(.a(dm_int_st2_27[3]), .b(dm_int_st2_27[4]), .cin(dm_int_st2_27[5]), .s(dm_int_st3_27[7]), .cout(dm_int_st3_28[1]));
	full_adder FA233(.a(dm_int_st2_27[6]), .b(dm_int_st2_27[7]), .cin(dm_int_st2_27[8]), .s(dm_int_st3_27[8]), .cout(dm_int_st3_28[2]));
	full_adder FA234(.a(dm_int_st2_27[9]), .b(dm_int_st2_27[10]), .cin(dm_int_st2_27[11]), .s(dm_int_st3_27[9]), .cout(dm_int_st3_28[3]));
	full_adder FA235(.a(dm_int_st2_27[12]), .b(dm_int_st2_27[13]), .cin(dm_int_st2_27[14]), .s(dm_int_st3_27[10]), .cout(dm_int_st3_28[4]));
	full_adder FA236(.a(dm_int_st2_27[15]), .b(dm_int_st2_27[16]), .cin(dm_int_st2_27[17]), .s(dm_int_st3_27[11]), .cout(dm_int_st3_28[5]));
	assign dm_int_st3_27[12] = dm_int_st2_27[18];
	// Bit 28
	full_adder FA237(.a(dm_int_st2_28[0]), .b(dm_int_st2_28[1]), .cin(dm_int_st2_28[2]), .s(dm_int_st3_28[6]), .cout(dm_int_st3_29[0]));
	full_adder FA238(.a(dm_int_st2_28[3]), .b(dm_int_st2_28[4]), .cin(dm_int_st2_28[5]), .s(dm_int_st3_28[7]), .cout(dm_int_st3_29[1]));
	full_adder FA239(.a(dm_int_st2_28[6]), .b(dm_int_st2_28[7]), .cin(dm_int_st2_28[8]), .s(dm_int_st3_28[8]), .cout(dm_int_st3_29[2]));
	full_adder FA240(.a(dm_int_st2_28[9]), .b(dm_int_st2_28[10]), .cin(dm_int_st2_28[11]), .s(dm_int_st3_28[9]), .cout(dm_int_st3_29[3]));
	full_adder FA241(.a(dm_int_st2_28[12]), .b(dm_int_st2_28[13]), .cin(dm_int_st2_28[14]), .s(dm_int_st3_28[10]), .cout(dm_int_st3_29[4]));
	full_adder FA242(.a(dm_int_st2_28[15]), .b(dm_int_st2_28[16]), .cin(dm_int_st2_28[17]), .s(dm_int_st3_28[11]), .cout(dm_int_st3_29[5]));
	assign dm_int_st3_28[12] = dm_int_st2_28[18];
	// Bit 29
	full_adder FA243(.a(dm_int_st2_29[0]), .b(dm_int_st2_29[1]), .cin(dm_int_st2_29[2]), .s(dm_int_st3_29[6]), .cout(dm_int_st3_30[0]));
	full_adder FA244(.a(dm_int_st2_29[3]), .b(dm_int_st2_29[4]), .cin(dm_int_st2_29[5]), .s(dm_int_st3_29[7]), .cout(dm_int_st3_30[1]));
	full_adder FA245(.a(dm_int_st2_29[6]), .b(dm_int_st2_29[7]), .cin(dm_int_st2_29[8]), .s(dm_int_st3_29[8]), .cout(dm_int_st3_30[2]));
	full_adder FA246(.a(dm_int_st2_29[9]), .b(dm_int_st2_29[10]), .cin(dm_int_st2_29[11]), .s(dm_int_st3_29[9]), .cout(dm_int_st3_30[3]));
	full_adder FA247(.a(dm_int_st2_29[12]), .b(dm_int_st2_29[13]), .cin(dm_int_st2_29[14]), .s(dm_int_st3_29[10]), .cout(dm_int_st3_30[4]));
	full_adder FA248(.a(dm_int_st2_29[15]), .b(dm_int_st2_29[16]), .cin(dm_int_st2_29[17]), .s(dm_int_st3_29[11]), .cout(dm_int_st3_30[5]));
	assign dm_int_st3_29[12] = dm_int_st2_29[18];
	// Bit 30
	full_adder FA249(.a(dm_int_st2_30[0]), .b(dm_int_st2_30[1]), .cin(dm_int_st2_30[2]), .s(dm_int_st3_30[6]), .cout(dm_int_st3_31[0]));
	full_adder FA250(.a(dm_int_st2_30[3]), .b(dm_int_st2_30[4]), .cin(dm_int_st2_30[5]), .s(dm_int_st3_30[7]), .cout(dm_int_st3_31[1]));
	full_adder FA251(.a(dm_int_st2_30[6]), .b(dm_int_st2_30[7]), .cin(dm_int_st2_30[8]), .s(dm_int_st3_30[8]), .cout(dm_int_st3_31[2]));
	full_adder FA252(.a(dm_int_st2_30[9]), .b(dm_int_st2_30[10]), .cin(dm_int_st2_30[11]), .s(dm_int_st3_30[9]), .cout(dm_int_st3_31[3]));
	full_adder FA253(.a(dm_int_st2_30[12]), .b(dm_int_st2_30[13]), .cin(dm_int_st2_30[14]), .s(dm_int_st3_30[10]), .cout(dm_int_st3_31[4]));
	full_adder FA254(.a(dm_int_st2_30[15]), .b(dm_int_st2_30[16]), .cin(dm_int_st2_30[17]), .s(dm_int_st3_30[11]), .cout(dm_int_st3_31[5]));
	assign dm_int_st3_30[12] = dm_int_st2_30[18];
	// Bit 31
	full_adder FA255(.a(dm_int_st2_31[0]), .b(dm_int_st2_31[1]), .cin(dm_int_st2_31[2]), .s(dm_int_st3_31[6]), .cout(dm_int_st3_32[0]));
	full_adder FA256(.a(dm_int_st2_31[3]), .b(dm_int_st2_31[4]), .cin(dm_int_st2_31[5]), .s(dm_int_st3_31[7]), .cout(dm_int_st3_32[1]));
	full_adder FA257(.a(dm_int_st2_31[6]), .b(dm_int_st2_31[7]), .cin(dm_int_st2_31[8]), .s(dm_int_st3_31[8]), .cout(dm_int_st3_32[2]));
	full_adder FA258(.a(dm_int_st2_31[9]), .b(dm_int_st2_31[10]), .cin(dm_int_st2_31[11]), .s(dm_int_st3_31[9]), .cout(dm_int_st3_32[3]));
	full_adder FA259(.a(dm_int_st2_31[12]), .b(dm_int_st2_31[13]), .cin(dm_int_st2_31[14]), .s(dm_int_st3_31[10]), .cout(dm_int_st3_32[4]));
	full_adder FA260(.a(dm_int_st2_31[15]), .b(dm_int_st2_31[16]), .cin(dm_int_st2_31[17]), .s(dm_int_st3_31[11]), .cout(dm_int_st3_32[5]));
	assign dm_int_st3_31[12] = dm_int_st2_31[18];
	// Bit 32
	full_adder FA261(.a(dm_int_st2_32[0]), .b(dm_int_st2_32[1]), .cin(dm_int_st2_32[2]), .s(dm_int_st3_32[6]), .cout(dm_int_st3_33[0]));
	full_adder FA262(.a(dm_int_st2_32[3]), .b(dm_int_st2_32[4]), .cin(dm_int_st2_32[5]), .s(dm_int_st3_32[7]), .cout(dm_int_st3_33[1]));
	full_adder FA263(.a(dm_int_st2_32[6]), .b(dm_int_st2_32[7]), .cin(dm_int_st2_32[8]), .s(dm_int_st3_32[8]), .cout(dm_int_st3_33[2]));
	full_adder FA264(.a(dm_int_st2_32[9]), .b(dm_int_st2_32[10]), .cin(dm_int_st2_32[11]), .s(dm_int_st3_32[9]), .cout(dm_int_st3_33[3]));
	full_adder FA265(.a(dm_int_st2_32[12]), .b(dm_int_st2_32[13]), .cin(dm_int_st2_32[14]), .s(dm_int_st3_32[10]), .cout(dm_int_st3_33[4]));
	full_adder FA266(.a(dm_int_st2_32[15]), .b(dm_int_st2_32[16]), .cin(dm_int_st2_32[17]), .s(dm_int_st3_32[11]), .cout(dm_int_st3_33[5]));
	assign dm_int_st3_32[12] = dm_int_st2_32[18];
	// Bit 33
	full_adder FA267(.a(dm_int_st2_33[0]), .b(dm_int_st2_33[1]), .cin(dm_int_st2_33[2]), .s(dm_int_st3_33[6]), .cout(dm_int_st3_34[0]));
	full_adder FA268(.a(dm_int_st2_33[3]), .b(dm_int_st2_33[4]), .cin(dm_int_st2_33[5]), .s(dm_int_st3_33[7]), .cout(dm_int_st3_34[1]));
	full_adder FA269(.a(dm_int_st2_33[6]), .b(dm_int_st2_33[7]), .cin(dm_int_st2_33[8]), .s(dm_int_st3_33[8]), .cout(dm_int_st3_34[2]));
	full_adder FA270(.a(dm_int_st2_33[9]), .b(dm_int_st2_33[10]), .cin(dm_int_st2_33[11]), .s(dm_int_st3_33[9]), .cout(dm_int_st3_34[3]));
	full_adder FA271(.a(dm_int_st2_33[12]), .b(dm_int_st2_33[13]), .cin(dm_int_st2_33[14]), .s(dm_int_st3_33[10]), .cout(dm_int_st3_34[4]));
	full_adder FA272(.a(dm_int_st2_33[15]), .b(dm_int_st2_33[16]), .cin(dm_int_st2_33[17]), .s(dm_int_st3_33[11]), .cout(dm_int_st3_34[5]));
	assign dm_int_st3_33[12] = dm_int_st2_33[18];
	// Bit 34
	full_adder FA273(.a(dm_int_st2_34[0]), .b(dm_int_st2_34[1]), .cin(dm_int_st2_34[2]), .s(dm_int_st3_34[6]), .cout(dm_int_st3_35[0]));
	full_adder FA274(.a(dm_int_st2_34[3]), .b(dm_int_st2_34[4]), .cin(dm_int_st2_34[5]), .s(dm_int_st3_34[7]), .cout(dm_int_st3_35[1]));
	full_adder FA275(.a(dm_int_st2_34[6]), .b(dm_int_st2_34[7]), .cin(dm_int_st2_34[8]), .s(dm_int_st3_34[8]), .cout(dm_int_st3_35[2]));
	full_adder FA276(.a(dm_int_st2_34[9]), .b(dm_int_st2_34[10]), .cin(dm_int_st2_34[11]), .s(dm_int_st3_34[9]), .cout(dm_int_st3_35[3]));
	full_adder FA277(.a(dm_int_st2_34[12]), .b(dm_int_st2_34[13]), .cin(dm_int_st2_34[14]), .s(dm_int_st3_34[10]), .cout(dm_int_st3_35[4]));
	full_adder FA278(.a(dm_int_st2_34[15]), .b(dm_int_st2_34[16]), .cin(dm_int_st2_34[17]), .s(dm_int_st3_34[11]), .cout(dm_int_st3_35[5]));
	assign dm_int_st3_34[12] = dm_int_st2_34[18];
	// Bit 35
	full_adder FA279(.a(dm_int_st2_35[0]), .b(dm_int_st2_35[1]), .cin(dm_int_st2_35[2]), .s(dm_int_st3_35[6]), .cout(dm_int_st3_36[0]));
	full_adder FA280(.a(dm_int_st2_35[3]), .b(dm_int_st2_35[4]), .cin(dm_int_st2_35[5]), .s(dm_int_st3_35[7]), .cout(dm_int_st3_36[1]));
	full_adder FA281(.a(dm_int_st2_35[6]), .b(dm_int_st2_35[7]), .cin(dm_int_st2_35[8]), .s(dm_int_st3_35[8]), .cout(dm_int_st3_36[2]));
	full_adder FA282(.a(dm_int_st2_35[9]), .b(dm_int_st2_35[10]), .cin(dm_int_st2_35[11]), .s(dm_int_st3_35[9]), .cout(dm_int_st3_36[3]));
	full_adder FA283(.a(dm_int_st2_35[12]), .b(dm_int_st2_35[13]), .cin(dm_int_st2_35[14]), .s(dm_int_st3_35[10]), .cout(dm_int_st3_36[4]));
	full_adder FA284(.a(dm_int_st2_35[15]), .b(dm_int_st2_35[16]), .cin(dm_int_st2_35[17]), .s(dm_int_st3_35[11]), .cout(dm_int_st3_36[5]));
	assign dm_int_st3_35[12] = dm_int_st2_35[18];
	// Bit 36
	full_adder FA285(.a(dm_int_st2_36[0]), .b(dm_int_st2_36[1]), .cin(dm_int_st2_36[2]), .s(dm_int_st3_36[6]), .cout(dm_int_st3_37[0]));
	full_adder FA286(.a(dm_int_st2_36[3]), .b(dm_int_st2_36[4]), .cin(dm_int_st2_36[5]), .s(dm_int_st3_36[7]), .cout(dm_int_st3_37[1]));
	full_adder FA287(.a(dm_int_st2_36[6]), .b(dm_int_st2_36[7]), .cin(dm_int_st2_36[8]), .s(dm_int_st3_36[8]), .cout(dm_int_st3_37[2]));
	full_adder FA288(.a(dm_int_st2_36[9]), .b(dm_int_st2_36[10]), .cin(dm_int_st2_36[11]), .s(dm_int_st3_36[9]), .cout(dm_int_st3_37[3]));
	full_adder FA289(.a(dm_int_st2_36[12]), .b(dm_int_st2_36[13]), .cin(dm_int_st2_36[14]), .s(dm_int_st3_36[10]), .cout(dm_int_st3_37[4]));
	full_adder FA290(.a(dm_int_st2_36[15]), .b(dm_int_st2_36[16]), .cin(dm_int_st2_36[17]), .s(dm_int_st3_36[11]), .cout(dm_int_st3_37[5]));
	assign dm_int_st3_36[12] = dm_int_st2_36[18];
	// Bit 37
	full_adder FA291(.a(dm_int_st2_37[0]), .b(dm_int_st2_37[1]), .cin(dm_int_st2_37[2]), .s(dm_int_st3_37[6]), .cout(dm_int_st3_38[0]));
	full_adder FA292(.a(dm_int_st2_37[3]), .b(dm_int_st2_37[4]), .cin(dm_int_st2_37[5]), .s(dm_int_st3_37[7]), .cout(dm_int_st3_38[1]));
	full_adder FA293(.a(dm_int_st2_37[6]), .b(dm_int_st2_37[7]), .cin(dm_int_st2_37[8]), .s(dm_int_st3_37[8]), .cout(dm_int_st3_38[2]));
	full_adder FA294(.a(dm_int_st2_37[9]), .b(dm_int_st2_37[10]), .cin(dm_int_st2_37[11]), .s(dm_int_st3_37[9]), .cout(dm_int_st3_38[3]));
	full_adder FA295(.a(dm_int_st2_37[12]), .b(dm_int_st2_37[13]), .cin(dm_int_st2_37[14]), .s(dm_int_st3_37[10]), .cout(dm_int_st3_38[4]));
	full_adder FA296(.a(dm_int_st2_37[15]), .b(dm_int_st2_37[16]), .cin(dm_int_st2_37[17]), .s(dm_int_st3_37[11]), .cout(dm_int_st3_38[5]));
	assign dm_int_st3_37[12] = dm_int_st2_37[18];
	// Bit 38
	full_adder FA297(.a(dm_int_st2_38[0]), .b(dm_int_st2_38[1]), .cin(dm_int_st2_38[2]), .s(dm_int_st3_38[6]), .cout(dm_int_st3_39[0]));
	full_adder FA298(.a(dm_int_st2_38[3]), .b(dm_int_st2_38[4]), .cin(dm_int_st2_38[5]), .s(dm_int_st3_38[7]), .cout(dm_int_st3_39[1]));
	full_adder FA299(.a(dm_int_st2_38[6]), .b(dm_int_st2_38[7]), .cin(dm_int_st2_38[8]), .s(dm_int_st3_38[8]), .cout(dm_int_st3_39[2]));
	full_adder FA300(.a(dm_int_st2_38[9]), .b(dm_int_st2_38[10]), .cin(dm_int_st2_38[11]), .s(dm_int_st3_38[9]), .cout(dm_int_st3_39[3]));
	full_adder FA301(.a(dm_int_st2_38[12]), .b(dm_int_st2_38[13]), .cin(dm_int_st2_38[14]), .s(dm_int_st3_38[10]), .cout(dm_int_st3_39[4]));
	full_adder FA302(.a(dm_int_st2_38[15]), .b(dm_int_st2_38[16]), .cin(dm_int_st2_38[17]), .s(dm_int_st3_38[11]), .cout(dm_int_st3_39[5]));
	assign dm_int_st3_38[12] = dm_int_st2_38[18];
	// Bit 39
	full_adder FA303(.a(dm_int_st2_39[0]), .b(dm_int_st2_39[1]), .cin(dm_int_st2_39[2]), .s(dm_int_st3_39[6]), .cout(dm_int_st3_40[0]));
	full_adder FA304(.a(dm_int_st2_39[3]), .b(dm_int_st2_39[4]), .cin(dm_int_st2_39[5]), .s(dm_int_st3_39[7]), .cout(dm_int_st3_40[1]));
	full_adder FA305(.a(dm_int_st2_39[6]), .b(dm_int_st2_39[7]), .cin(dm_int_st2_39[8]), .s(dm_int_st3_39[8]), .cout(dm_int_st3_40[2]));
	full_adder FA306(.a(dm_int_st2_39[9]), .b(dm_int_st2_39[10]), .cin(dm_int_st2_39[11]), .s(dm_int_st3_39[9]), .cout(dm_int_st3_40[3]));
	full_adder FA307(.a(dm_int_st2_39[12]), .b(dm_int_st2_39[13]), .cin(dm_int_st2_39[14]), .s(dm_int_st3_39[10]), .cout(dm_int_st3_40[4]));
	full_adder FA308(.a(dm_int_st2_39[15]), .b(dm_int_st2_39[16]), .cin(dm_int_st2_39[17]), .s(dm_int_st3_39[11]), .cout(dm_int_st3_40[5]));
	assign dm_int_st3_39[12] = dm_int_st2_39[18];
	// Bit 40
	full_adder FA309(.a(dm_int_st2_40[0]), .b(dm_int_st2_40[1]), .cin(dm_int_st2_40[2]), .s(dm_int_st3_40[6]), .cout(dm_int_st3_41[0]));
	full_adder FA310(.a(dm_int_st2_40[3]), .b(dm_int_st2_40[4]), .cin(dm_int_st2_40[5]), .s(dm_int_st3_40[7]), .cout(dm_int_st3_41[1]));
	full_adder FA311(.a(dm_int_st2_40[6]), .b(dm_int_st2_40[7]), .cin(dm_int_st2_40[8]), .s(dm_int_st3_40[8]), .cout(dm_int_st3_41[2]));
	full_adder FA312(.a(dm_int_st2_40[9]), .b(dm_int_st2_40[10]), .cin(dm_int_st2_40[11]), .s(dm_int_st3_40[9]), .cout(dm_int_st3_41[3]));
	full_adder FA313(.a(dm_int_st2_40[12]), .b(dm_int_st2_40[13]), .cin(dm_int_st2_40[14]), .s(dm_int_st3_40[10]), .cout(dm_int_st3_41[4]));
	full_adder FA314(.a(dm_int_st2_40[15]), .b(dm_int_st2_40[16]), .cin(dm_int_st2_40[17]), .s(dm_int_st3_40[11]), .cout(dm_int_st3_41[5]));
	assign dm_int_st3_40[12] = dm_int_st2_40[18];
	// Bit 41
	full_adder FA315(.a(dm_int_st2_41[0]), .b(dm_int_st2_41[1]), .cin(dm_int_st2_41[2]), .s(dm_int_st3_41[6]), .cout(dm_int_st3_42[0]));
	full_adder FA316(.a(dm_int_st2_41[3]), .b(dm_int_st2_41[4]), .cin(dm_int_st2_41[5]), .s(dm_int_st3_41[7]), .cout(dm_int_st3_42[1]));
	full_adder FA317(.a(dm_int_st2_41[6]), .b(dm_int_st2_41[7]), .cin(dm_int_st2_41[8]), .s(dm_int_st3_41[8]), .cout(dm_int_st3_42[2]));
	full_adder FA318(.a(dm_int_st2_41[9]), .b(dm_int_st2_41[10]), .cin(dm_int_st2_41[11]), .s(dm_int_st3_41[9]), .cout(dm_int_st3_42[3]));
	full_adder FA319(.a(dm_int_st2_41[12]), .b(dm_int_st2_41[13]), .cin(dm_int_st2_41[14]), .s(dm_int_st3_41[10]), .cout(dm_int_st3_42[4]));
	full_adder FA320(.a(dm_int_st2_41[15]), .b(dm_int_st2_41[16]), .cin(dm_int_st2_41[17]), .s(dm_int_st3_41[11]), .cout(dm_int_st3_42[5]));
	assign dm_int_st3_41[12] = dm_int_st2_41[18];
	// Bit 42
	full_adder FA321(.a(dm_int_st2_42[0]), .b(dm_int_st2_42[1]), .cin(dm_int_st2_42[2]), .s(dm_int_st3_42[6]), .cout(dm_int_st3_43[0]));
	full_adder FA322(.a(dm_int_st2_42[3]), .b(dm_int_st2_42[4]), .cin(dm_int_st2_42[5]), .s(dm_int_st3_42[7]), .cout(dm_int_st3_43[1]));
	full_adder FA323(.a(dm_int_st2_42[6]), .b(dm_int_st2_42[7]), .cin(dm_int_st2_42[8]), .s(dm_int_st3_42[8]), .cout(dm_int_st3_43[2]));
	full_adder FA324(.a(dm_int_st2_42[9]), .b(dm_int_st2_42[10]), .cin(dm_int_st2_42[11]), .s(dm_int_st3_42[9]), .cout(dm_int_st3_43[3]));
	full_adder FA325(.a(dm_int_st2_42[12]), .b(dm_int_st2_42[13]), .cin(dm_int_st2_42[14]), .s(dm_int_st3_42[10]), .cout(dm_int_st3_43[4]));
	full_adder FA326(.a(dm_int_st2_42[15]), .b(dm_int_st2_42[16]), .cin(dm_int_st2_42[17]), .s(dm_int_st3_42[11]), .cout(dm_int_st3_43[5]));
	assign dm_int_st3_42[12] = dm_int_st2_42[18];
	// Bit 43
	full_adder FA327(.a(dm_int_st2_43[0]), .b(dm_int_st2_43[1]), .cin(dm_int_st2_43[2]), .s(dm_int_st3_43[6]), .cout(dm_int_st3_44[0]));
	full_adder FA328(.a(dm_int_st2_43[3]), .b(dm_int_st2_43[4]), .cin(dm_int_st2_43[5]), .s(dm_int_st3_43[7]), .cout(dm_int_st3_44[1]));
	full_adder FA329(.a(dm_int_st2_43[6]), .b(dm_int_st2_43[7]), .cin(dm_int_st2_43[8]), .s(dm_int_st3_43[8]), .cout(dm_int_st3_44[2]));
	full_adder FA330(.a(dm_int_st2_43[9]), .b(dm_int_st2_43[10]), .cin(dm_int_st2_43[11]), .s(dm_int_st3_43[9]), .cout(dm_int_st3_44[3]));
	full_adder FA331(.a(dm_int_st2_43[12]), .b(dm_int_st2_43[13]), .cin(dm_int_st2_43[14]), .s(dm_int_st3_43[10]), .cout(dm_int_st3_44[4]));
	full_adder FA332(.a(dm_int_st2_43[15]), .b(dm_int_st2_43[16]), .cin(dm_int_st2_43[17]), .s(dm_int_st3_43[11]), .cout(dm_int_st3_44[5]));
	assign dm_int_st3_43[12] = dm_int_st2_43[18];
	// Bit 44
	full_adder FA333(.a(dm_int_st2_44[0]), .b(dm_int_st2_44[1]), .cin(dm_int_st2_44[2]), .s(dm_int_st3_44[6]), .cout(dm_int_st3_45[0]));
	full_adder FA334(.a(dm_int_st2_44[3]), .b(dm_int_st2_44[4]), .cin(dm_int_st2_44[5]), .s(dm_int_st3_44[7]), .cout(dm_int_st3_45[1]));
	full_adder FA335(.a(dm_int_st2_44[6]), .b(dm_int_st2_44[7]), .cin(dm_int_st2_44[8]), .s(dm_int_st3_44[8]), .cout(dm_int_st3_45[2]));
	full_adder FA336(.a(dm_int_st2_44[9]), .b(dm_int_st2_44[10]), .cin(dm_int_st2_44[11]), .s(dm_int_st3_44[9]), .cout(dm_int_st3_45[3]));
	full_adder FA337(.a(dm_int_st2_44[12]), .b(dm_int_st2_44[13]), .cin(dm_int_st2_44[14]), .s(dm_int_st3_44[10]), .cout(dm_int_st3_45[4]));
	full_adder FA338(.a(dm_int_st2_44[15]), .b(dm_int_st2_44[16]), .cin(dm_int_st2_44[17]), .s(dm_int_st3_44[11]), .cout(dm_int_st3_45[5]));
	assign dm_int_st3_44[12] = dm_int_st2_44[18];
	// Bit 45
	full_adder FA339(.a(dm_int_st2_45[0]), .b(dm_int_st2_45[1]), .cin(dm_int_st2_45[2]), .s(dm_int_st3_45[6]), .cout(dm_int_st3_46[0]));
	full_adder FA340(.a(dm_int_st2_45[3]), .b(dm_int_st2_45[4]), .cin(dm_int_st2_45[5]), .s(dm_int_st3_45[7]), .cout(dm_int_st3_46[1]));
	full_adder FA341(.a(dm_int_st2_45[6]), .b(dm_int_st2_45[7]), .cin(dm_int_st2_45[8]), .s(dm_int_st3_45[8]), .cout(dm_int_st3_46[2]));
	full_adder FA342(.a(dm_int_st2_45[9]), .b(dm_int_st2_45[10]), .cin(dm_int_st2_45[11]), .s(dm_int_st3_45[9]), .cout(dm_int_st3_46[3]));
	full_adder FA343(.a(dm_int_st2_45[12]), .b(dm_int_st2_45[13]), .cin(dm_int_st2_45[14]), .s(dm_int_st3_45[10]), .cout(dm_int_st3_46[4]));
	full_adder FA344(.a(dm_int_st2_45[15]), .b(dm_int_st2_45[16]), .cin(dm_int_st2_45[17]), .s(dm_int_st3_45[11]), .cout(dm_int_st3_46[5]));
	assign dm_int_st3_45[12] = dm_int_st2_45[18];
	// Bit 46
	full_adder FA345(.a(dm_int_st2_46[0]), .b(dm_int_st2_46[1]), .cin(dm_int_st2_46[2]), .s(dm_int_st3_46[6]), .cout(dm_int_st3_47[0]));
	full_adder FA346(.a(dm_int_st2_46[3]), .b(dm_int_st2_46[4]), .cin(dm_int_st2_46[5]), .s(dm_int_st3_46[7]), .cout(dm_int_st3_47[1]));
	full_adder FA347(.a(dm_int_st2_46[6]), .b(dm_int_st2_46[7]), .cin(dm_int_st2_46[8]), .s(dm_int_st3_46[8]), .cout(dm_int_st3_47[2]));
	full_adder FA348(.a(dm_int_st2_46[9]), .b(dm_int_st2_46[10]), .cin(dm_int_st2_46[11]), .s(dm_int_st3_46[9]), .cout(dm_int_st3_47[3]));
	full_adder FA349(.a(dm_int_st2_46[12]), .b(dm_int_st2_46[13]), .cin(dm_int_st2_46[14]), .s(dm_int_st3_46[10]), .cout(dm_int_st3_47[4]));
	assign dm_int_st3_46[11] = dm_int_st2_46[15];
	assign dm_int_st3_46[12] = dm_int_st2_46[16];
	// Bit 47
	full_adder FA350(.a(dm_int_st2_47[0]), .b(dm_int_st2_47[1]), .cin(dm_int_st2_47[2]), .s(dm_int_st3_47[5]), .cout(dm_int_st3_48[0]));
	full_adder FA351(.a(dm_int_st2_47[3]), .b(dm_int_st2_47[4]), .cin(dm_int_st2_47[5]), .s(dm_int_st3_47[6]), .cout(dm_int_st3_48[1]));
	full_adder FA352(.a(dm_int_st2_47[6]), .b(dm_int_st2_47[7]), .cin(dm_int_st2_47[8]), .s(dm_int_st3_47[7]), .cout(dm_int_st3_48[2]));
	full_adder FA353(.a(dm_int_st2_47[9]), .b(dm_int_st2_47[10]), .cin(dm_int_st2_47[11]), .s(dm_int_st3_47[8]), .cout(dm_int_st3_48[3]));
	assign dm_int_st3_47[9] = dm_int_st2_47[12];
	assign dm_int_st3_47[10] = dm_int_st2_47[13];
	assign dm_int_st3_47[11] = dm_int_st2_47[14];
	assign dm_int_st3_47[12] = dm_int_st2_47[15];
	// Bit 48
	full_adder FA354(.a(dm_int_st2_48[0]), .b(dm_int_st2_48[1]), .cin(dm_int_st2_48[2]), .s(dm_int_st3_48[4]), .cout(dm_int_st3_49[0]));
	full_adder FA355(.a(dm_int_st2_48[3]), .b(dm_int_st2_48[4]), .cin(dm_int_st2_48[5]), .s(dm_int_st3_48[5]), .cout(dm_int_st3_49[1]));
	full_adder FA356(.a(dm_int_st2_48[6]), .b(dm_int_st2_48[7]), .cin(dm_int_st2_48[8]), .s(dm_int_st3_48[6]), .cout(dm_int_st3_49[2]));
	assign dm_int_st3_48[7] = dm_int_st2_48[9];
	assign dm_int_st3_48[8] = dm_int_st2_48[10];
	assign dm_int_st3_48[9] = dm_int_st2_48[11];
	assign dm_int_st3_48[10] = dm_int_st2_48[12];
	assign dm_int_st3_48[11] = dm_int_st2_48[13];
	assign dm_int_st3_48[12] = dm_int_st2_48[14];
	// Bit 49
	full_adder FA357(.a(dm_int_st2_49[0]), .b(dm_int_st2_49[1]), .cin(dm_int_st2_49[2]), .s(dm_int_st3_49[3]), .cout(dm_int_st3_50[0]));
	full_adder FA358(.a(dm_int_st2_49[3]), .b(dm_int_st2_49[4]), .cin(dm_int_st2_49[5]), .s(dm_int_st3_49[4]), .cout(dm_int_st3_50[1]));
	assign dm_int_st3_49[5] = dm_int_st2_49[6];
	assign dm_int_st3_49[6] = dm_int_st2_49[7];
	assign dm_int_st3_49[7] = dm_int_st2_49[8];
	assign dm_int_st3_49[8] = dm_int_st2_49[9];
	assign dm_int_st3_49[9] = dm_int_st2_49[10];
	assign dm_int_st3_49[10] = dm_int_st2_49[11];
	assign dm_int_st3_49[11] = dm_int_st2_49[12];
	assign dm_int_st3_49[12] = dm_int_st2_49[13];
	// Bit 50
	full_adder FA359(.a(dm_int_st2_50[0]), .b(dm_int_st2_50[1]), .cin(dm_int_st2_50[2]), .s(dm_int_st3_50[2]), .cout(dm_int_st3_51[0]));
	assign dm_int_st3_50[3] = dm_int_st2_50[3];
	assign dm_int_st3_50[4] = dm_int_st2_50[4];
	assign dm_int_st3_50[5] = dm_int_st2_50[5];
	assign dm_int_st3_50[6] = dm_int_st2_50[6];
	assign dm_int_st3_50[7] = dm_int_st2_50[7];
	assign dm_int_st3_50[8] = dm_int_st2_50[8];
	assign dm_int_st3_50[9] = dm_int_st2_50[9];
	assign dm_int_st3_50[10] = dm_int_st2_50[10];
	assign dm_int_st3_50[11] = dm_int_st2_50[11];
	assign dm_int_st3_50[12] = dm_int_st2_50[12];
	// Bit 51
	assign dm_int_st3_51[1] = dm_int_st2_51[0];
	assign dm_int_st3_51[2] = dm_int_st2_51[1];
	assign dm_int_st3_51[3] = dm_int_st2_51[2];
	assign dm_int_st3_51[4] = dm_int_st2_51[3];
	assign dm_int_st3_51[5] = dm_int_st2_51[4];
	assign dm_int_st3_51[6] = dm_int_st2_51[5];
	assign dm_int_st3_51[7] = dm_int_st2_51[6];
	assign dm_int_st3_51[8] = dm_int_st2_51[7];
	assign dm_int_st3_51[9] = dm_int_st2_51[8];
	assign dm_int_st3_51[10] = dm_int_st2_51[9];
	assign dm_int_st3_51[11] = dm_int_st2_51[10];
	assign dm_int_st3_51[12] = dm_int_st2_51[11];
	// Bit 52
	assign dm_int_st3_52[0] = dm_int_st2_52[0];
	assign dm_int_st3_52[1] = dm_int_st2_52[1];
	assign dm_int_st3_52[2] = dm_int_st2_52[2];
	assign dm_int_st3_52[3] = dm_int_st2_52[3];
	assign dm_int_st3_52[4] = dm_int_st2_52[4];
	assign dm_int_st3_52[5] = dm_int_st2_52[5];
	assign dm_int_st3_52[6] = dm_int_st2_52[6];
	assign dm_int_st3_52[7] = dm_int_st2_52[7];
	assign dm_int_st3_52[8] = dm_int_st2_52[8];
	assign dm_int_st3_52[9] = dm_int_st2_52[9];
	assign dm_int_st3_52[10] = dm_int_st2_52[10];
	// Bit 53
	assign dm_int_st3_53[0] = dm_int_st2_53[0];
	assign dm_int_st3_53[1] = dm_int_st2_53[1];
	assign dm_int_st3_53[2] = dm_int_st2_53[2];
	assign dm_int_st3_53[3] = dm_int_st2_53[3];
	assign dm_int_st3_53[4] = dm_int_st2_53[4];
	assign dm_int_st3_53[5] = dm_int_st2_53[5];
	assign dm_int_st3_53[6] = dm_int_st2_53[6];
	assign dm_int_st3_53[7] = dm_int_st2_53[7];
	assign dm_int_st3_53[8] = dm_int_st2_53[8];
	assign dm_int_st3_53[9] = dm_int_st2_53[9];
	// Bit 54
	assign dm_int_st3_54[0] = dm_int_st2_54[0];
	assign dm_int_st3_54[1] = dm_int_st2_54[1];
	assign dm_int_st3_54[2] = dm_int_st2_54[2];
	assign dm_int_st3_54[3] = dm_int_st2_54[3];
	assign dm_int_st3_54[4] = dm_int_st2_54[4];
	assign dm_int_st3_54[5] = dm_int_st2_54[5];
	assign dm_int_st3_54[6] = dm_int_st2_54[6];
	assign dm_int_st3_54[7] = dm_int_st2_54[7];
	assign dm_int_st3_54[8] = dm_int_st2_54[8];
	// Bit 55
	assign dm_int_st3_55[0] = dm_int_st2_55[0];
	assign dm_int_st3_55[1] = dm_int_st2_55[1];
	assign dm_int_st3_55[2] = dm_int_st2_55[2];
	assign dm_int_st3_55[3] = dm_int_st2_55[3];
	assign dm_int_st3_55[4] = dm_int_st2_55[4];
	assign dm_int_st3_55[5] = dm_int_st2_55[5];
	assign dm_int_st3_55[6] = dm_int_st2_55[6];
	assign dm_int_st3_55[7] = dm_int_st2_55[7];
	// Bit 56
	assign dm_int_st3_56[0] = dm_int_st2_56[0];
	assign dm_int_st3_56[1] = dm_int_st2_56[1];
	assign dm_int_st3_56[2] = dm_int_st2_56[2];
	assign dm_int_st3_56[3] = dm_int_st2_56[3];
	assign dm_int_st3_56[4] = dm_int_st2_56[4];
	assign dm_int_st3_56[5] = dm_int_st2_56[5];
	assign dm_int_st3_56[6] = dm_int_st2_56[6];
	// Bit 57
	assign dm_int_st3_57[0] = dm_int_st2_57[0];
	assign dm_int_st3_57[1] = dm_int_st2_57[1];
	assign dm_int_st3_57[2] = dm_int_st2_57[2];
	assign dm_int_st3_57[3] = dm_int_st2_57[3];
	assign dm_int_st3_57[4] = dm_int_st2_57[4];
	assign dm_int_st3_57[5] = dm_int_st2_57[5];
	// Bit 58
	assign dm_int_st3_58[0] = dm_int_st2_58[0];
	assign dm_int_st3_58[1] = dm_int_st2_58[1];
	assign dm_int_st3_58[2] = dm_int_st2_58[2];
	assign dm_int_st3_58[3] = dm_int_st2_58[3];
	assign dm_int_st3_58[4] = dm_int_st2_58[4];
	// Bit 59
	assign dm_int_st3_59[0] = dm_int_st2_59[0];
	assign dm_int_st3_59[1] = dm_int_st2_59[1];
	assign dm_int_st3_59[2] = dm_int_st2_59[2];
	assign dm_int_st3_59[3] = dm_int_st2_59[3];
	// Bit 60
	assign dm_int_st3_60[0] = dm_int_st2_60[0];
	assign dm_int_st3_60[1] = dm_int_st2_60[1];
	assign dm_int_st3_60[2] = dm_int_st2_60[2];
	// Bit 61
	assign dm_int_st3_61[0] = dm_int_st2_61[0];
	assign dm_int_st3_61[1] = dm_int_st2_61[1];
	// Bit 62
	assign dm_int_st3_62[0] = dm_int_st2_62[0];

	//// Stage 4 ////
	wire [0:0] dm_int_st4_0;
	wire [1:0] dm_int_st4_1;
	wire [2:0] dm_int_st4_2;
	wire [3:0] dm_int_st4_3;
	wire [4:0] dm_int_st4_4;
	wire [5:0] dm_int_st4_5;
	wire [6:0] dm_int_st4_6;
	wire [7:0] dm_int_st4_7;
	wire [8:0] dm_int_st4_8;
	wire [8:0] dm_int_st4_9;
	wire [8:0] dm_int_st4_10;
	wire [8:0] dm_int_st4_11;
	wire [8:0] dm_int_st4_12;
	wire [8:0] dm_int_st4_13;
	wire [8:0] dm_int_st4_14;
	wire [8:0] dm_int_st4_15;
	wire [8:0] dm_int_st4_16;
	wire [8:0] dm_int_st4_17;
	wire [8:0] dm_int_st4_18;
	wire [8:0] dm_int_st4_19;
	wire [8:0] dm_int_st4_20;
	wire [8:0] dm_int_st4_21;
	wire [8:0] dm_int_st4_22;
	wire [8:0] dm_int_st4_23;
	wire [8:0] dm_int_st4_24;
	wire [8:0] dm_int_st4_25;
	wire [8:0] dm_int_st4_26;
	wire [8:0] dm_int_st4_27;
	wire [8:0] dm_int_st4_28;
	wire [8:0] dm_int_st4_29;
	wire [8:0] dm_int_st4_30;
	wire [8:0] dm_int_st4_31;
	wire [8:0] dm_int_st4_32;
	wire [8:0] dm_int_st4_33;
	wire [8:0] dm_int_st4_34;
	wire [8:0] dm_int_st4_35;
	wire [8:0] dm_int_st4_36;
	wire [8:0] dm_int_st4_37;
	wire [8:0] dm_int_st4_38;
	wire [8:0] dm_int_st4_39;
	wire [8:0] dm_int_st4_40;
	wire [8:0] dm_int_st4_41;
	wire [8:0] dm_int_st4_42;
	wire [8:0] dm_int_st4_43;
	wire [8:0] dm_int_st4_44;
	wire [8:0] dm_int_st4_45;
	wire [8:0] dm_int_st4_46;
	wire [8:0] dm_int_st4_47;
	wire [8:0] dm_int_st4_48;
	wire [8:0] dm_int_st4_49;
	wire [8:0] dm_int_st4_50;
	wire [8:0] dm_int_st4_51;
	wire [8:0] dm_int_st4_52;
	wire [8:0] dm_int_st4_53;
	wire [8:0] dm_int_st4_54;
	wire [8:0] dm_int_st4_55;
	wire [6:0] dm_int_st4_56;
	wire [5:0] dm_int_st4_57;
	wire [4:0] dm_int_st4_58;
	wire [3:0] dm_int_st4_59;
	wire [2:0] dm_int_st4_60;
	wire [1:0] dm_int_st4_61;
	wire [0:0] dm_int_st4_62;

	// Bit 0
	assign dm_int_st4_0[0] = dm_int_st3_0[0];
	// Bit 1
	assign dm_int_st4_1[0] = dm_int_st3_1[0];
	assign dm_int_st4_1[1] = dm_int_st3_1[1];
	// Bit 2
	assign dm_int_st4_2[0] = dm_int_st3_2[0];
	assign dm_int_st4_2[1] = dm_int_st3_2[1];
	assign dm_int_st4_2[2] = dm_int_st3_2[2];
	// Bit 3
	assign dm_int_st4_3[0] = dm_int_st3_3[0];
	assign dm_int_st4_3[1] = dm_int_st3_3[1];
	assign dm_int_st4_3[2] = dm_int_st3_3[2];
	assign dm_int_st4_3[3] = dm_int_st3_3[3];
	// Bit 4
	assign dm_int_st4_4[0] = dm_int_st3_4[0];
	assign dm_int_st4_4[1] = dm_int_st3_4[1];
	assign dm_int_st4_4[2] = dm_int_st3_4[2];
	assign dm_int_st4_4[3] = dm_int_st3_4[3];
	assign dm_int_st4_4[4] = dm_int_st3_4[4];
	// Bit 5
	assign dm_int_st4_5[0] = dm_int_st3_5[0];
	assign dm_int_st4_5[1] = dm_int_st3_5[1];
	assign dm_int_st4_5[2] = dm_int_st3_5[2];
	assign dm_int_st4_5[3] = dm_int_st3_5[3];
	assign dm_int_st4_5[4] = dm_int_st3_5[4];
	assign dm_int_st4_5[5] = dm_int_st3_5[5];
	// Bit 6
	assign dm_int_st4_6[0] = dm_int_st3_6[0];
	assign dm_int_st4_6[1] = dm_int_st3_6[1];
	assign dm_int_st4_6[2] = dm_int_st3_6[2];
	assign dm_int_st4_6[3] = dm_int_st3_6[3];
	assign dm_int_st4_6[4] = dm_int_st3_6[4];
	assign dm_int_st4_6[5] = dm_int_st3_6[5];
	assign dm_int_st4_6[6] = dm_int_st3_6[6];
	// Bit 7
	assign dm_int_st4_7[0] = dm_int_st3_7[0];
	assign dm_int_st4_7[1] = dm_int_st3_7[1];
	assign dm_int_st4_7[2] = dm_int_st3_7[2];
	assign dm_int_st4_7[3] = dm_int_st3_7[3];
	assign dm_int_st4_7[4] = dm_int_st3_7[4];
	assign dm_int_st4_7[5] = dm_int_st3_7[5];
	assign dm_int_st4_7[6] = dm_int_st3_7[6];
	assign dm_int_st4_7[7] = dm_int_st3_7[7];
	// Bit 8
	assign dm_int_st4_8[0] = dm_int_st3_8[0];
	assign dm_int_st4_8[1] = dm_int_st3_8[1];
	assign dm_int_st4_8[2] = dm_int_st3_8[2];
	assign dm_int_st4_8[3] = dm_int_st3_8[3];
	assign dm_int_st4_8[4] = dm_int_st3_8[4];
	assign dm_int_st4_8[5] = dm_int_st3_8[5];
	assign dm_int_st4_8[6] = dm_int_st3_8[6];
	assign dm_int_st4_8[7] = dm_int_st3_8[7];
	assign dm_int_st4_8[8] = dm_int_st3_8[8];
	// Bit 9
	half_adder HA20(.a(dm_int_st3_9[0]), .b(dm_int_st3_9[1]), .s(dm_int_st4_9[0]), .cout(dm_int_st4_10[0]));
	assign dm_int_st4_9[1] = dm_int_st3_9[2];
	assign dm_int_st4_9[2] = dm_int_st3_9[3];
	assign dm_int_st4_9[3] = dm_int_st3_9[4];
	assign dm_int_st4_9[4] = dm_int_st3_9[5];
	assign dm_int_st4_9[5] = dm_int_st3_9[6];
	assign dm_int_st4_9[6] = dm_int_st3_9[7];
	assign dm_int_st4_9[7] = dm_int_st3_9[8];
	assign dm_int_st4_9[8] = dm_int_st3_9[9];
	// Bit 10
	full_adder FA360(.a(dm_int_st3_10[0]), .b(dm_int_st3_10[1]), .cin(dm_int_st3_10[2]), .s(dm_int_st4_10[1]), .cout(dm_int_st4_11[0]));
	half_adder HA21(.a(dm_int_st3_10[3]), .b(dm_int_st3_10[4]), .s(dm_int_st4_10[2]), .cout(dm_int_st4_11[1]));
	assign dm_int_st4_10[3] = dm_int_st3_10[5];
	assign dm_int_st4_10[4] = dm_int_st3_10[6];
	assign dm_int_st4_10[5] = dm_int_st3_10[7];
	assign dm_int_st4_10[6] = dm_int_st3_10[8];
	assign dm_int_st4_10[7] = dm_int_st3_10[9];
	assign dm_int_st4_10[8] = dm_int_st3_10[10];
	// Bit 11
	full_adder FA361(.a(dm_int_st3_11[0]), .b(dm_int_st3_11[1]), .cin(dm_int_st3_11[2]), .s(dm_int_st4_11[2]), .cout(dm_int_st4_12[0]));
	full_adder FA362(.a(dm_int_st3_11[3]), .b(dm_int_st3_11[4]), .cin(dm_int_st3_11[5]), .s(dm_int_st4_11[3]), .cout(dm_int_st4_12[1]));
	half_adder HA22(.a(dm_int_st3_11[6]), .b(dm_int_st3_11[7]), .s(dm_int_st4_11[4]), .cout(dm_int_st4_12[2]));
	assign dm_int_st4_11[5] = dm_int_st3_11[8];
	assign dm_int_st4_11[6] = dm_int_st3_11[9];
	assign dm_int_st4_11[7] = dm_int_st3_11[10];
	assign dm_int_st4_11[8] = dm_int_st3_11[11];
	// Bit 12
	full_adder FA363(.a(dm_int_st3_12[0]), .b(dm_int_st3_12[1]), .cin(dm_int_st3_12[2]), .s(dm_int_st4_12[3]), .cout(dm_int_st4_13[0]));
	full_adder FA364(.a(dm_int_st3_12[3]), .b(dm_int_st3_12[4]), .cin(dm_int_st3_12[5]), .s(dm_int_st4_12[4]), .cout(dm_int_st4_13[1]));
	full_adder FA365(.a(dm_int_st3_12[6]), .b(dm_int_st3_12[7]), .cin(dm_int_st3_12[8]), .s(dm_int_st4_12[5]), .cout(dm_int_st4_13[2]));
	half_adder HA23(.a(dm_int_st3_12[9]), .b(dm_int_st3_12[10]), .s(dm_int_st4_12[6]), .cout(dm_int_st4_13[3]));
	assign dm_int_st4_12[7] = dm_int_st3_12[11];
	assign dm_int_st4_12[8] = dm_int_st3_12[12];
	// Bit 13
	full_adder FA366(.a(dm_int_st3_13[0]), .b(dm_int_st3_13[1]), .cin(dm_int_st3_13[2]), .s(dm_int_st4_13[4]), .cout(dm_int_st4_14[0]));
	full_adder FA367(.a(dm_int_st3_13[3]), .b(dm_int_st3_13[4]), .cin(dm_int_st3_13[5]), .s(dm_int_st4_13[5]), .cout(dm_int_st4_14[1]));
	full_adder FA368(.a(dm_int_st3_13[6]), .b(dm_int_st3_13[7]), .cin(dm_int_st3_13[8]), .s(dm_int_st4_13[6]), .cout(dm_int_st4_14[2]));
	full_adder FA369(.a(dm_int_st3_13[9]), .b(dm_int_st3_13[10]), .cin(dm_int_st3_13[11]), .s(dm_int_st4_13[7]), .cout(dm_int_st4_14[3]));
	assign dm_int_st4_13[8] = dm_int_st3_13[12];
	// Bit 14
	full_adder FA370(.a(dm_int_st3_14[0]), .b(dm_int_st3_14[1]), .cin(dm_int_st3_14[2]), .s(dm_int_st4_14[4]), .cout(dm_int_st4_15[0]));
	full_adder FA371(.a(dm_int_st3_14[3]), .b(dm_int_st3_14[4]), .cin(dm_int_st3_14[5]), .s(dm_int_st4_14[5]), .cout(dm_int_st4_15[1]));
	full_adder FA372(.a(dm_int_st3_14[6]), .b(dm_int_st3_14[7]), .cin(dm_int_st3_14[8]), .s(dm_int_st4_14[6]), .cout(dm_int_st4_15[2]));
	full_adder FA373(.a(dm_int_st3_14[9]), .b(dm_int_st3_14[10]), .cin(dm_int_st3_14[11]), .s(dm_int_st4_14[7]), .cout(dm_int_st4_15[3]));
	assign dm_int_st4_14[8] = dm_int_st3_14[12];
	// Bit 15
	full_adder FA374(.a(dm_int_st3_15[0]), .b(dm_int_st3_15[1]), .cin(dm_int_st3_15[2]), .s(dm_int_st4_15[4]), .cout(dm_int_st4_16[0]));
	full_adder FA375(.a(dm_int_st3_15[3]), .b(dm_int_st3_15[4]), .cin(dm_int_st3_15[5]), .s(dm_int_st4_15[5]), .cout(dm_int_st4_16[1]));
	full_adder FA376(.a(dm_int_st3_15[6]), .b(dm_int_st3_15[7]), .cin(dm_int_st3_15[8]), .s(dm_int_st4_15[6]), .cout(dm_int_st4_16[2]));
	full_adder FA377(.a(dm_int_st3_15[9]), .b(dm_int_st3_15[10]), .cin(dm_int_st3_15[11]), .s(dm_int_st4_15[7]), .cout(dm_int_st4_16[3]));
	assign dm_int_st4_15[8] = dm_int_st3_15[12];
	// Bit 16
	full_adder FA378(.a(dm_int_st3_16[0]), .b(dm_int_st3_16[1]), .cin(dm_int_st3_16[2]), .s(dm_int_st4_16[4]), .cout(dm_int_st4_17[0]));
	full_adder FA379(.a(dm_int_st3_16[3]), .b(dm_int_st3_16[4]), .cin(dm_int_st3_16[5]), .s(dm_int_st4_16[5]), .cout(dm_int_st4_17[1]));
	full_adder FA380(.a(dm_int_st3_16[6]), .b(dm_int_st3_16[7]), .cin(dm_int_st3_16[8]), .s(dm_int_st4_16[6]), .cout(dm_int_st4_17[2]));
	full_adder FA381(.a(dm_int_st3_16[9]), .b(dm_int_st3_16[10]), .cin(dm_int_st3_16[11]), .s(dm_int_st4_16[7]), .cout(dm_int_st4_17[3]));
	assign dm_int_st4_16[8] = dm_int_st3_16[12];
	// Bit 17
	full_adder FA382(.a(dm_int_st3_17[0]), .b(dm_int_st3_17[1]), .cin(dm_int_st3_17[2]), .s(dm_int_st4_17[4]), .cout(dm_int_st4_18[0]));
	full_adder FA383(.a(dm_int_st3_17[3]), .b(dm_int_st3_17[4]), .cin(dm_int_st3_17[5]), .s(dm_int_st4_17[5]), .cout(dm_int_st4_18[1]));
	full_adder FA384(.a(dm_int_st3_17[6]), .b(dm_int_st3_17[7]), .cin(dm_int_st3_17[8]), .s(dm_int_st4_17[6]), .cout(dm_int_st4_18[2]));
	full_adder FA385(.a(dm_int_st3_17[9]), .b(dm_int_st3_17[10]), .cin(dm_int_st3_17[11]), .s(dm_int_st4_17[7]), .cout(dm_int_st4_18[3]));
	assign dm_int_st4_17[8] = dm_int_st3_17[12];
	// Bit 18
	full_adder FA386(.a(dm_int_st3_18[0]), .b(dm_int_st3_18[1]), .cin(dm_int_st3_18[2]), .s(dm_int_st4_18[4]), .cout(dm_int_st4_19[0]));
	full_adder FA387(.a(dm_int_st3_18[3]), .b(dm_int_st3_18[4]), .cin(dm_int_st3_18[5]), .s(dm_int_st4_18[5]), .cout(dm_int_st4_19[1]));
	full_adder FA388(.a(dm_int_st3_18[6]), .b(dm_int_st3_18[7]), .cin(dm_int_st3_18[8]), .s(dm_int_st4_18[6]), .cout(dm_int_st4_19[2]));
	full_adder FA389(.a(dm_int_st3_18[9]), .b(dm_int_st3_18[10]), .cin(dm_int_st3_18[11]), .s(dm_int_st4_18[7]), .cout(dm_int_st4_19[3]));
	assign dm_int_st4_18[8] = dm_int_st3_18[12];
	// Bit 19
	full_adder FA390(.a(dm_int_st3_19[0]), .b(dm_int_st3_19[1]), .cin(dm_int_st3_19[2]), .s(dm_int_st4_19[4]), .cout(dm_int_st4_20[0]));
	full_adder FA391(.a(dm_int_st3_19[3]), .b(dm_int_st3_19[4]), .cin(dm_int_st3_19[5]), .s(dm_int_st4_19[5]), .cout(dm_int_st4_20[1]));
	full_adder FA392(.a(dm_int_st3_19[6]), .b(dm_int_st3_19[7]), .cin(dm_int_st3_19[8]), .s(dm_int_st4_19[6]), .cout(dm_int_st4_20[2]));
	full_adder FA393(.a(dm_int_st3_19[9]), .b(dm_int_st3_19[10]), .cin(dm_int_st3_19[11]), .s(dm_int_st4_19[7]), .cout(dm_int_st4_20[3]));
	assign dm_int_st4_19[8] = dm_int_st3_19[12];
	// Bit 20
	full_adder FA394(.a(dm_int_st3_20[0]), .b(dm_int_st3_20[1]), .cin(dm_int_st3_20[2]), .s(dm_int_st4_20[4]), .cout(dm_int_st4_21[0]));
	full_adder FA395(.a(dm_int_st3_20[3]), .b(dm_int_st3_20[4]), .cin(dm_int_st3_20[5]), .s(dm_int_st4_20[5]), .cout(dm_int_st4_21[1]));
	full_adder FA396(.a(dm_int_st3_20[6]), .b(dm_int_st3_20[7]), .cin(dm_int_st3_20[8]), .s(dm_int_st4_20[6]), .cout(dm_int_st4_21[2]));
	full_adder FA397(.a(dm_int_st3_20[9]), .b(dm_int_st3_20[10]), .cin(dm_int_st3_20[11]), .s(dm_int_st4_20[7]), .cout(dm_int_st4_21[3]));
	assign dm_int_st4_20[8] = dm_int_st3_20[12];
	// Bit 21
	full_adder FA398(.a(dm_int_st3_21[0]), .b(dm_int_st3_21[1]), .cin(dm_int_st3_21[2]), .s(dm_int_st4_21[4]), .cout(dm_int_st4_22[0]));
	full_adder FA399(.a(dm_int_st3_21[3]), .b(dm_int_st3_21[4]), .cin(dm_int_st3_21[5]), .s(dm_int_st4_21[5]), .cout(dm_int_st4_22[1]));
	full_adder FA400(.a(dm_int_st3_21[6]), .b(dm_int_st3_21[7]), .cin(dm_int_st3_21[8]), .s(dm_int_st4_21[6]), .cout(dm_int_st4_22[2]));
	full_adder FA401(.a(dm_int_st3_21[9]), .b(dm_int_st3_21[10]), .cin(dm_int_st3_21[11]), .s(dm_int_st4_21[7]), .cout(dm_int_st4_22[3]));
	assign dm_int_st4_21[8] = dm_int_st3_21[12];
	// Bit 22
	full_adder FA402(.a(dm_int_st3_22[0]), .b(dm_int_st3_22[1]), .cin(dm_int_st3_22[2]), .s(dm_int_st4_22[4]), .cout(dm_int_st4_23[0]));
	full_adder FA403(.a(dm_int_st3_22[3]), .b(dm_int_st3_22[4]), .cin(dm_int_st3_22[5]), .s(dm_int_st4_22[5]), .cout(dm_int_st4_23[1]));
	full_adder FA404(.a(dm_int_st3_22[6]), .b(dm_int_st3_22[7]), .cin(dm_int_st3_22[8]), .s(dm_int_st4_22[6]), .cout(dm_int_st4_23[2]));
	full_adder FA405(.a(dm_int_st3_22[9]), .b(dm_int_st3_22[10]), .cin(dm_int_st3_22[11]), .s(dm_int_st4_22[7]), .cout(dm_int_st4_23[3]));
	assign dm_int_st4_22[8] = dm_int_st3_22[12];
	// Bit 23
	full_adder FA406(.a(dm_int_st3_23[0]), .b(dm_int_st3_23[1]), .cin(dm_int_st3_23[2]), .s(dm_int_st4_23[4]), .cout(dm_int_st4_24[0]));
	full_adder FA407(.a(dm_int_st3_23[3]), .b(dm_int_st3_23[4]), .cin(dm_int_st3_23[5]), .s(dm_int_st4_23[5]), .cout(dm_int_st4_24[1]));
	full_adder FA408(.a(dm_int_st3_23[6]), .b(dm_int_st3_23[7]), .cin(dm_int_st3_23[8]), .s(dm_int_st4_23[6]), .cout(dm_int_st4_24[2]));
	full_adder FA409(.a(dm_int_st3_23[9]), .b(dm_int_st3_23[10]), .cin(dm_int_st3_23[11]), .s(dm_int_st4_23[7]), .cout(dm_int_st4_24[3]));
	assign dm_int_st4_23[8] = dm_int_st3_23[12];
	// Bit 24
	full_adder FA410(.a(dm_int_st3_24[0]), .b(dm_int_st3_24[1]), .cin(dm_int_st3_24[2]), .s(dm_int_st4_24[4]), .cout(dm_int_st4_25[0]));
	full_adder FA411(.a(dm_int_st3_24[3]), .b(dm_int_st3_24[4]), .cin(dm_int_st3_24[5]), .s(dm_int_st4_24[5]), .cout(dm_int_st4_25[1]));
	full_adder FA412(.a(dm_int_st3_24[6]), .b(dm_int_st3_24[7]), .cin(dm_int_st3_24[8]), .s(dm_int_st4_24[6]), .cout(dm_int_st4_25[2]));
	full_adder FA413(.a(dm_int_st3_24[9]), .b(dm_int_st3_24[10]), .cin(dm_int_st3_24[11]), .s(dm_int_st4_24[7]), .cout(dm_int_st4_25[3]));
	assign dm_int_st4_24[8] = dm_int_st3_24[12];
	// Bit 25
	full_adder FA414(.a(dm_int_st3_25[0]), .b(dm_int_st3_25[1]), .cin(dm_int_st3_25[2]), .s(dm_int_st4_25[4]), .cout(dm_int_st4_26[0]));
	full_adder FA415(.a(dm_int_st3_25[3]), .b(dm_int_st3_25[4]), .cin(dm_int_st3_25[5]), .s(dm_int_st4_25[5]), .cout(dm_int_st4_26[1]));
	full_adder FA416(.a(dm_int_st3_25[6]), .b(dm_int_st3_25[7]), .cin(dm_int_st3_25[8]), .s(dm_int_st4_25[6]), .cout(dm_int_st4_26[2]));
	full_adder FA417(.a(dm_int_st3_25[9]), .b(dm_int_st3_25[10]), .cin(dm_int_st3_25[11]), .s(dm_int_st4_25[7]), .cout(dm_int_st4_26[3]));
	assign dm_int_st4_25[8] = dm_int_st3_25[12];
	// Bit 26
	full_adder FA418(.a(dm_int_st3_26[0]), .b(dm_int_st3_26[1]), .cin(dm_int_st3_26[2]), .s(dm_int_st4_26[4]), .cout(dm_int_st4_27[0]));
	full_adder FA419(.a(dm_int_st3_26[3]), .b(dm_int_st3_26[4]), .cin(dm_int_st3_26[5]), .s(dm_int_st4_26[5]), .cout(dm_int_st4_27[1]));
	full_adder FA420(.a(dm_int_st3_26[6]), .b(dm_int_st3_26[7]), .cin(dm_int_st3_26[8]), .s(dm_int_st4_26[6]), .cout(dm_int_st4_27[2]));
	full_adder FA421(.a(dm_int_st3_26[9]), .b(dm_int_st3_26[10]), .cin(dm_int_st3_26[11]), .s(dm_int_st4_26[7]), .cout(dm_int_st4_27[3]));
	assign dm_int_st4_26[8] = dm_int_st3_26[12];
	// Bit 27
	full_adder FA422(.a(dm_int_st3_27[0]), .b(dm_int_st3_27[1]), .cin(dm_int_st3_27[2]), .s(dm_int_st4_27[4]), .cout(dm_int_st4_28[0]));
	full_adder FA423(.a(dm_int_st3_27[3]), .b(dm_int_st3_27[4]), .cin(dm_int_st3_27[5]), .s(dm_int_st4_27[5]), .cout(dm_int_st4_28[1]));
	full_adder FA424(.a(dm_int_st3_27[6]), .b(dm_int_st3_27[7]), .cin(dm_int_st3_27[8]), .s(dm_int_st4_27[6]), .cout(dm_int_st4_28[2]));
	full_adder FA425(.a(dm_int_st3_27[9]), .b(dm_int_st3_27[10]), .cin(dm_int_st3_27[11]), .s(dm_int_st4_27[7]), .cout(dm_int_st4_28[3]));
	assign dm_int_st4_27[8] = dm_int_st3_27[12];
	// Bit 28
	full_adder FA426(.a(dm_int_st3_28[0]), .b(dm_int_st3_28[1]), .cin(dm_int_st3_28[2]), .s(dm_int_st4_28[4]), .cout(dm_int_st4_29[0]));
	full_adder FA427(.a(dm_int_st3_28[3]), .b(dm_int_st3_28[4]), .cin(dm_int_st3_28[5]), .s(dm_int_st4_28[5]), .cout(dm_int_st4_29[1]));
	full_adder FA428(.a(dm_int_st3_28[6]), .b(dm_int_st3_28[7]), .cin(dm_int_st3_28[8]), .s(dm_int_st4_28[6]), .cout(dm_int_st4_29[2]));
	full_adder FA429(.a(dm_int_st3_28[9]), .b(dm_int_st3_28[10]), .cin(dm_int_st3_28[11]), .s(dm_int_st4_28[7]), .cout(dm_int_st4_29[3]));
	assign dm_int_st4_28[8] = dm_int_st3_28[12];
	// Bit 29
	full_adder FA430(.a(dm_int_st3_29[0]), .b(dm_int_st3_29[1]), .cin(dm_int_st3_29[2]), .s(dm_int_st4_29[4]), .cout(dm_int_st4_30[0]));
	full_adder FA431(.a(dm_int_st3_29[3]), .b(dm_int_st3_29[4]), .cin(dm_int_st3_29[5]), .s(dm_int_st4_29[5]), .cout(dm_int_st4_30[1]));
	full_adder FA432(.a(dm_int_st3_29[6]), .b(dm_int_st3_29[7]), .cin(dm_int_st3_29[8]), .s(dm_int_st4_29[6]), .cout(dm_int_st4_30[2]));
	full_adder FA433(.a(dm_int_st3_29[9]), .b(dm_int_st3_29[10]), .cin(dm_int_st3_29[11]), .s(dm_int_st4_29[7]), .cout(dm_int_st4_30[3]));
	assign dm_int_st4_29[8] = dm_int_st3_29[12];
	// Bit 30
	full_adder FA434(.a(dm_int_st3_30[0]), .b(dm_int_st3_30[1]), .cin(dm_int_st3_30[2]), .s(dm_int_st4_30[4]), .cout(dm_int_st4_31[0]));
	full_adder FA435(.a(dm_int_st3_30[3]), .b(dm_int_st3_30[4]), .cin(dm_int_st3_30[5]), .s(dm_int_st4_30[5]), .cout(dm_int_st4_31[1]));
	full_adder FA436(.a(dm_int_st3_30[6]), .b(dm_int_st3_30[7]), .cin(dm_int_st3_30[8]), .s(dm_int_st4_30[6]), .cout(dm_int_st4_31[2]));
	full_adder FA437(.a(dm_int_st3_30[9]), .b(dm_int_st3_30[10]), .cin(dm_int_st3_30[11]), .s(dm_int_st4_30[7]), .cout(dm_int_st4_31[3]));
	assign dm_int_st4_30[8] = dm_int_st3_30[12];
	// Bit 31
	full_adder FA438(.a(dm_int_st3_31[0]), .b(dm_int_st3_31[1]), .cin(dm_int_st3_31[2]), .s(dm_int_st4_31[4]), .cout(dm_int_st4_32[0]));
	full_adder FA439(.a(dm_int_st3_31[3]), .b(dm_int_st3_31[4]), .cin(dm_int_st3_31[5]), .s(dm_int_st4_31[5]), .cout(dm_int_st4_32[1]));
	full_adder FA440(.a(dm_int_st3_31[6]), .b(dm_int_st3_31[7]), .cin(dm_int_st3_31[8]), .s(dm_int_st4_31[6]), .cout(dm_int_st4_32[2]));
	full_adder FA441(.a(dm_int_st3_31[9]), .b(dm_int_st3_31[10]), .cin(dm_int_st3_31[11]), .s(dm_int_st4_31[7]), .cout(dm_int_st4_32[3]));
	assign dm_int_st4_31[8] = dm_int_st3_31[12];
	// Bit 32
	full_adder FA442(.a(dm_int_st3_32[0]), .b(dm_int_st3_32[1]), .cin(dm_int_st3_32[2]), .s(dm_int_st4_32[4]), .cout(dm_int_st4_33[0]));
	full_adder FA443(.a(dm_int_st3_32[3]), .b(dm_int_st3_32[4]), .cin(dm_int_st3_32[5]), .s(dm_int_st4_32[5]), .cout(dm_int_st4_33[1]));
	full_adder FA444(.a(dm_int_st3_32[6]), .b(dm_int_st3_32[7]), .cin(dm_int_st3_32[8]), .s(dm_int_st4_32[6]), .cout(dm_int_st4_33[2]));
	full_adder FA445(.a(dm_int_st3_32[9]), .b(dm_int_st3_32[10]), .cin(dm_int_st3_32[11]), .s(dm_int_st4_32[7]), .cout(dm_int_st4_33[3]));
	assign dm_int_st4_32[8] = dm_int_st3_32[12];
	// Bit 33
	full_adder FA446(.a(dm_int_st3_33[0]), .b(dm_int_st3_33[1]), .cin(dm_int_st3_33[2]), .s(dm_int_st4_33[4]), .cout(dm_int_st4_34[0]));
	full_adder FA447(.a(dm_int_st3_33[3]), .b(dm_int_st3_33[4]), .cin(dm_int_st3_33[5]), .s(dm_int_st4_33[5]), .cout(dm_int_st4_34[1]));
	full_adder FA448(.a(dm_int_st3_33[6]), .b(dm_int_st3_33[7]), .cin(dm_int_st3_33[8]), .s(dm_int_st4_33[6]), .cout(dm_int_st4_34[2]));
	full_adder FA449(.a(dm_int_st3_33[9]), .b(dm_int_st3_33[10]), .cin(dm_int_st3_33[11]), .s(dm_int_st4_33[7]), .cout(dm_int_st4_34[3]));
	assign dm_int_st4_33[8] = dm_int_st3_33[12];
	// Bit 34
	full_adder FA450(.a(dm_int_st3_34[0]), .b(dm_int_st3_34[1]), .cin(dm_int_st3_34[2]), .s(dm_int_st4_34[4]), .cout(dm_int_st4_35[0]));
	full_adder FA451(.a(dm_int_st3_34[3]), .b(dm_int_st3_34[4]), .cin(dm_int_st3_34[5]), .s(dm_int_st4_34[5]), .cout(dm_int_st4_35[1]));
	full_adder FA452(.a(dm_int_st3_34[6]), .b(dm_int_st3_34[7]), .cin(dm_int_st3_34[8]), .s(dm_int_st4_34[6]), .cout(dm_int_st4_35[2]));
	full_adder FA453(.a(dm_int_st3_34[9]), .b(dm_int_st3_34[10]), .cin(dm_int_st3_34[11]), .s(dm_int_st4_34[7]), .cout(dm_int_st4_35[3]));
	assign dm_int_st4_34[8] = dm_int_st3_34[12];
	// Bit 35
	full_adder FA454(.a(dm_int_st3_35[0]), .b(dm_int_st3_35[1]), .cin(dm_int_st3_35[2]), .s(dm_int_st4_35[4]), .cout(dm_int_st4_36[0]));
	full_adder FA455(.a(dm_int_st3_35[3]), .b(dm_int_st3_35[4]), .cin(dm_int_st3_35[5]), .s(dm_int_st4_35[5]), .cout(dm_int_st4_36[1]));
	full_adder FA456(.a(dm_int_st3_35[6]), .b(dm_int_st3_35[7]), .cin(dm_int_st3_35[8]), .s(dm_int_st4_35[6]), .cout(dm_int_st4_36[2]));
	full_adder FA457(.a(dm_int_st3_35[9]), .b(dm_int_st3_35[10]), .cin(dm_int_st3_35[11]), .s(dm_int_st4_35[7]), .cout(dm_int_st4_36[3]));
	assign dm_int_st4_35[8] = dm_int_st3_35[12];
	// Bit 36
	full_adder FA458(.a(dm_int_st3_36[0]), .b(dm_int_st3_36[1]), .cin(dm_int_st3_36[2]), .s(dm_int_st4_36[4]), .cout(dm_int_st4_37[0]));
	full_adder FA459(.a(dm_int_st3_36[3]), .b(dm_int_st3_36[4]), .cin(dm_int_st3_36[5]), .s(dm_int_st4_36[5]), .cout(dm_int_st4_37[1]));
	full_adder FA460(.a(dm_int_st3_36[6]), .b(dm_int_st3_36[7]), .cin(dm_int_st3_36[8]), .s(dm_int_st4_36[6]), .cout(dm_int_st4_37[2]));
	full_adder FA461(.a(dm_int_st3_36[9]), .b(dm_int_st3_36[10]), .cin(dm_int_st3_36[11]), .s(dm_int_st4_36[7]), .cout(dm_int_st4_37[3]));
	assign dm_int_st4_36[8] = dm_int_st3_36[12];
	// Bit 37
	full_adder FA462(.a(dm_int_st3_37[0]), .b(dm_int_st3_37[1]), .cin(dm_int_st3_37[2]), .s(dm_int_st4_37[4]), .cout(dm_int_st4_38[0]));
	full_adder FA463(.a(dm_int_st3_37[3]), .b(dm_int_st3_37[4]), .cin(dm_int_st3_37[5]), .s(dm_int_st4_37[5]), .cout(dm_int_st4_38[1]));
	full_adder FA464(.a(dm_int_st3_37[6]), .b(dm_int_st3_37[7]), .cin(dm_int_st3_37[8]), .s(dm_int_st4_37[6]), .cout(dm_int_st4_38[2]));
	full_adder FA465(.a(dm_int_st3_37[9]), .b(dm_int_st3_37[10]), .cin(dm_int_st3_37[11]), .s(dm_int_st4_37[7]), .cout(dm_int_st4_38[3]));
	assign dm_int_st4_37[8] = dm_int_st3_37[12];
	// Bit 38
	full_adder FA466(.a(dm_int_st3_38[0]), .b(dm_int_st3_38[1]), .cin(dm_int_st3_38[2]), .s(dm_int_st4_38[4]), .cout(dm_int_st4_39[0]));
	full_adder FA467(.a(dm_int_st3_38[3]), .b(dm_int_st3_38[4]), .cin(dm_int_st3_38[5]), .s(dm_int_st4_38[5]), .cout(dm_int_st4_39[1]));
	full_adder FA468(.a(dm_int_st3_38[6]), .b(dm_int_st3_38[7]), .cin(dm_int_st3_38[8]), .s(dm_int_st4_38[6]), .cout(dm_int_st4_39[2]));
	full_adder FA469(.a(dm_int_st3_38[9]), .b(dm_int_st3_38[10]), .cin(dm_int_st3_38[11]), .s(dm_int_st4_38[7]), .cout(dm_int_st4_39[3]));
	assign dm_int_st4_38[8] = dm_int_st3_38[12];
	// Bit 39
	full_adder FA470(.a(dm_int_st3_39[0]), .b(dm_int_st3_39[1]), .cin(dm_int_st3_39[2]), .s(dm_int_st4_39[4]), .cout(dm_int_st4_40[0]));
	full_adder FA471(.a(dm_int_st3_39[3]), .b(dm_int_st3_39[4]), .cin(dm_int_st3_39[5]), .s(dm_int_st4_39[5]), .cout(dm_int_st4_40[1]));
	full_adder FA472(.a(dm_int_st3_39[6]), .b(dm_int_st3_39[7]), .cin(dm_int_st3_39[8]), .s(dm_int_st4_39[6]), .cout(dm_int_st4_40[2]));
	full_adder FA473(.a(dm_int_st3_39[9]), .b(dm_int_st3_39[10]), .cin(dm_int_st3_39[11]), .s(dm_int_st4_39[7]), .cout(dm_int_st4_40[3]));
	assign dm_int_st4_39[8] = dm_int_st3_39[12];
	// Bit 40
	full_adder FA474(.a(dm_int_st3_40[0]), .b(dm_int_st3_40[1]), .cin(dm_int_st3_40[2]), .s(dm_int_st4_40[4]), .cout(dm_int_st4_41[0]));
	full_adder FA475(.a(dm_int_st3_40[3]), .b(dm_int_st3_40[4]), .cin(dm_int_st3_40[5]), .s(dm_int_st4_40[5]), .cout(dm_int_st4_41[1]));
	full_adder FA476(.a(dm_int_st3_40[6]), .b(dm_int_st3_40[7]), .cin(dm_int_st3_40[8]), .s(dm_int_st4_40[6]), .cout(dm_int_st4_41[2]));
	full_adder FA477(.a(dm_int_st3_40[9]), .b(dm_int_st3_40[10]), .cin(dm_int_st3_40[11]), .s(dm_int_st4_40[7]), .cout(dm_int_st4_41[3]));
	assign dm_int_st4_40[8] = dm_int_st3_40[12];
	// Bit 41
	full_adder FA478(.a(dm_int_st3_41[0]), .b(dm_int_st3_41[1]), .cin(dm_int_st3_41[2]), .s(dm_int_st4_41[4]), .cout(dm_int_st4_42[0]));
	full_adder FA479(.a(dm_int_st3_41[3]), .b(dm_int_st3_41[4]), .cin(dm_int_st3_41[5]), .s(dm_int_st4_41[5]), .cout(dm_int_st4_42[1]));
	full_adder FA480(.a(dm_int_st3_41[6]), .b(dm_int_st3_41[7]), .cin(dm_int_st3_41[8]), .s(dm_int_st4_41[6]), .cout(dm_int_st4_42[2]));
	full_adder FA481(.a(dm_int_st3_41[9]), .b(dm_int_st3_41[10]), .cin(dm_int_st3_41[11]), .s(dm_int_st4_41[7]), .cout(dm_int_st4_42[3]));
	assign dm_int_st4_41[8] = dm_int_st3_41[12];
	// Bit 42
	full_adder FA482(.a(dm_int_st3_42[0]), .b(dm_int_st3_42[1]), .cin(dm_int_st3_42[2]), .s(dm_int_st4_42[4]), .cout(dm_int_st4_43[0]));
	full_adder FA483(.a(dm_int_st3_42[3]), .b(dm_int_st3_42[4]), .cin(dm_int_st3_42[5]), .s(dm_int_st4_42[5]), .cout(dm_int_st4_43[1]));
	full_adder FA484(.a(dm_int_st3_42[6]), .b(dm_int_st3_42[7]), .cin(dm_int_st3_42[8]), .s(dm_int_st4_42[6]), .cout(dm_int_st4_43[2]));
	full_adder FA485(.a(dm_int_st3_42[9]), .b(dm_int_st3_42[10]), .cin(dm_int_st3_42[11]), .s(dm_int_st4_42[7]), .cout(dm_int_st4_43[3]));
	assign dm_int_st4_42[8] = dm_int_st3_42[12];
	// Bit 43
	full_adder FA486(.a(dm_int_st3_43[0]), .b(dm_int_st3_43[1]), .cin(dm_int_st3_43[2]), .s(dm_int_st4_43[4]), .cout(dm_int_st4_44[0]));
	full_adder FA487(.a(dm_int_st3_43[3]), .b(dm_int_st3_43[4]), .cin(dm_int_st3_43[5]), .s(dm_int_st4_43[5]), .cout(dm_int_st4_44[1]));
	full_adder FA488(.a(dm_int_st3_43[6]), .b(dm_int_st3_43[7]), .cin(dm_int_st3_43[8]), .s(dm_int_st4_43[6]), .cout(dm_int_st4_44[2]));
	full_adder FA489(.a(dm_int_st3_43[9]), .b(dm_int_st3_43[10]), .cin(dm_int_st3_43[11]), .s(dm_int_st4_43[7]), .cout(dm_int_st4_44[3]));
	assign dm_int_st4_43[8] = dm_int_st3_43[12];
	// Bit 44
	full_adder FA490(.a(dm_int_st3_44[0]), .b(dm_int_st3_44[1]), .cin(dm_int_st3_44[2]), .s(dm_int_st4_44[4]), .cout(dm_int_st4_45[0]));
	full_adder FA491(.a(dm_int_st3_44[3]), .b(dm_int_st3_44[4]), .cin(dm_int_st3_44[5]), .s(dm_int_st4_44[5]), .cout(dm_int_st4_45[1]));
	full_adder FA492(.a(dm_int_st3_44[6]), .b(dm_int_st3_44[7]), .cin(dm_int_st3_44[8]), .s(dm_int_st4_44[6]), .cout(dm_int_st4_45[2]));
	full_adder FA493(.a(dm_int_st3_44[9]), .b(dm_int_st3_44[10]), .cin(dm_int_st3_44[11]), .s(dm_int_st4_44[7]), .cout(dm_int_st4_45[3]));
	assign dm_int_st4_44[8] = dm_int_st3_44[12];
	// Bit 45
	full_adder FA494(.a(dm_int_st3_45[0]), .b(dm_int_st3_45[1]), .cin(dm_int_st3_45[2]), .s(dm_int_st4_45[4]), .cout(dm_int_st4_46[0]));
	full_adder FA495(.a(dm_int_st3_45[3]), .b(dm_int_st3_45[4]), .cin(dm_int_st3_45[5]), .s(dm_int_st4_45[5]), .cout(dm_int_st4_46[1]));
	full_adder FA496(.a(dm_int_st3_45[6]), .b(dm_int_st3_45[7]), .cin(dm_int_st3_45[8]), .s(dm_int_st4_45[6]), .cout(dm_int_st4_46[2]));
	full_adder FA497(.a(dm_int_st3_45[9]), .b(dm_int_st3_45[10]), .cin(dm_int_st3_45[11]), .s(dm_int_st4_45[7]), .cout(dm_int_st4_46[3]));
	assign dm_int_st4_45[8] = dm_int_st3_45[12];
	// Bit 46
	full_adder FA498(.a(dm_int_st3_46[0]), .b(dm_int_st3_46[1]), .cin(dm_int_st3_46[2]), .s(dm_int_st4_46[4]), .cout(dm_int_st4_47[0]));
	full_adder FA499(.a(dm_int_st3_46[3]), .b(dm_int_st3_46[4]), .cin(dm_int_st3_46[5]), .s(dm_int_st4_46[5]), .cout(dm_int_st4_47[1]));
	full_adder FA500(.a(dm_int_st3_46[6]), .b(dm_int_st3_46[7]), .cin(dm_int_st3_46[8]), .s(dm_int_st4_46[6]), .cout(dm_int_st4_47[2]));
	full_adder FA501(.a(dm_int_st3_46[9]), .b(dm_int_st3_46[10]), .cin(dm_int_st3_46[11]), .s(dm_int_st4_46[7]), .cout(dm_int_st4_47[3]));
	assign dm_int_st4_46[8] = dm_int_st3_46[12];
	// Bit 47
	full_adder FA502(.a(dm_int_st3_47[0]), .b(dm_int_st3_47[1]), .cin(dm_int_st3_47[2]), .s(dm_int_st4_47[4]), .cout(dm_int_st4_48[0]));
	full_adder FA503(.a(dm_int_st3_47[3]), .b(dm_int_st3_47[4]), .cin(dm_int_st3_47[5]), .s(dm_int_st4_47[5]), .cout(dm_int_st4_48[1]));
	full_adder FA504(.a(dm_int_st3_47[6]), .b(dm_int_st3_47[7]), .cin(dm_int_st3_47[8]), .s(dm_int_st4_47[6]), .cout(dm_int_st4_48[2]));
	full_adder FA505(.a(dm_int_st3_47[9]), .b(dm_int_st3_47[10]), .cin(dm_int_st3_47[11]), .s(dm_int_st4_47[7]), .cout(dm_int_st4_48[3]));
	assign dm_int_st4_47[8] = dm_int_st3_47[12];
	// Bit 48
	full_adder FA506(.a(dm_int_st3_48[0]), .b(dm_int_st3_48[1]), .cin(dm_int_st3_48[2]), .s(dm_int_st4_48[4]), .cout(dm_int_st4_49[0]));
	full_adder FA507(.a(dm_int_st3_48[3]), .b(dm_int_st3_48[4]), .cin(dm_int_st3_48[5]), .s(dm_int_st4_48[5]), .cout(dm_int_st4_49[1]));
	full_adder FA508(.a(dm_int_st3_48[6]), .b(dm_int_st3_48[7]), .cin(dm_int_st3_48[8]), .s(dm_int_st4_48[6]), .cout(dm_int_st4_49[2]));
	full_adder FA509(.a(dm_int_st3_48[9]), .b(dm_int_st3_48[10]), .cin(dm_int_st3_48[11]), .s(dm_int_st4_48[7]), .cout(dm_int_st4_49[3]));
	assign dm_int_st4_48[8] = dm_int_st3_48[12];
	// Bit 49
	full_adder FA510(.a(dm_int_st3_49[0]), .b(dm_int_st3_49[1]), .cin(dm_int_st3_49[2]), .s(dm_int_st4_49[4]), .cout(dm_int_st4_50[0]));
	full_adder FA511(.a(dm_int_st3_49[3]), .b(dm_int_st3_49[4]), .cin(dm_int_st3_49[5]), .s(dm_int_st4_49[5]), .cout(dm_int_st4_50[1]));
	full_adder FA512(.a(dm_int_st3_49[6]), .b(dm_int_st3_49[7]), .cin(dm_int_st3_49[8]), .s(dm_int_st4_49[6]), .cout(dm_int_st4_50[2]));
	full_adder FA513(.a(dm_int_st3_49[9]), .b(dm_int_st3_49[10]), .cin(dm_int_st3_49[11]), .s(dm_int_st4_49[7]), .cout(dm_int_st4_50[3]));
	assign dm_int_st4_49[8] = dm_int_st3_49[12];
	// Bit 50
	full_adder FA514(.a(dm_int_st3_50[0]), .b(dm_int_st3_50[1]), .cin(dm_int_st3_50[2]), .s(dm_int_st4_50[4]), .cout(dm_int_st4_51[0]));
	full_adder FA515(.a(dm_int_st3_50[3]), .b(dm_int_st3_50[4]), .cin(dm_int_st3_50[5]), .s(dm_int_st4_50[5]), .cout(dm_int_st4_51[1]));
	full_adder FA516(.a(dm_int_st3_50[6]), .b(dm_int_st3_50[7]), .cin(dm_int_st3_50[8]), .s(dm_int_st4_50[6]), .cout(dm_int_st4_51[2]));
	full_adder FA517(.a(dm_int_st3_50[9]), .b(dm_int_st3_50[10]), .cin(dm_int_st3_50[11]), .s(dm_int_st4_50[7]), .cout(dm_int_st4_51[3]));
	assign dm_int_st4_50[8] = dm_int_st3_50[12];
	// Bit 51
	full_adder FA518(.a(dm_int_st3_51[0]), .b(dm_int_st3_51[1]), .cin(dm_int_st3_51[2]), .s(dm_int_st4_51[4]), .cout(dm_int_st4_52[0]));
	full_adder FA519(.a(dm_int_st3_51[3]), .b(dm_int_st3_51[4]), .cin(dm_int_st3_51[5]), .s(dm_int_st4_51[5]), .cout(dm_int_st4_52[1]));
	full_adder FA520(.a(dm_int_st3_51[6]), .b(dm_int_st3_51[7]), .cin(dm_int_st3_51[8]), .s(dm_int_st4_51[6]), .cout(dm_int_st4_52[2]));
	full_adder FA521(.a(dm_int_st3_51[9]), .b(dm_int_st3_51[10]), .cin(dm_int_st3_51[11]), .s(dm_int_st4_51[7]), .cout(dm_int_st4_52[3]));
	assign dm_int_st4_51[8] = dm_int_st3_51[12];
	// Bit 52
	full_adder FA522(.a(dm_int_st3_52[0]), .b(dm_int_st3_52[1]), .cin(dm_int_st3_52[2]), .s(dm_int_st4_52[4]), .cout(dm_int_st4_53[0]));
	full_adder FA523(.a(dm_int_st3_52[3]), .b(dm_int_st3_52[4]), .cin(dm_int_st3_52[5]), .s(dm_int_st4_52[5]), .cout(dm_int_st4_53[1]));
	full_adder FA524(.a(dm_int_st3_52[6]), .b(dm_int_st3_52[7]), .cin(dm_int_st3_52[8]), .s(dm_int_st4_52[6]), .cout(dm_int_st4_53[2]));
	assign dm_int_st4_52[7] = dm_int_st3_52[9];
	assign dm_int_st4_52[8] = dm_int_st3_52[10];
	// Bit 53
	full_adder FA525(.a(dm_int_st3_53[0]), .b(dm_int_st3_53[1]), .cin(dm_int_st3_53[2]), .s(dm_int_st4_53[3]), .cout(dm_int_st4_54[0]));
	full_adder FA526(.a(dm_int_st3_53[3]), .b(dm_int_st3_53[4]), .cin(dm_int_st3_53[5]), .s(dm_int_st4_53[4]), .cout(dm_int_st4_54[1]));
	assign dm_int_st4_53[5] = dm_int_st3_53[6];
	assign dm_int_st4_53[6] = dm_int_st3_53[7];
	assign dm_int_st4_53[7] = dm_int_st3_53[8];
	assign dm_int_st4_53[8] = dm_int_st3_53[9];
	// Bit 54
	full_adder FA527(.a(dm_int_st3_54[0]), .b(dm_int_st3_54[1]), .cin(dm_int_st3_54[2]), .s(dm_int_st4_54[2]), .cout(dm_int_st4_55[0]));
	assign dm_int_st4_54[3] = dm_int_st3_54[3];
	assign dm_int_st4_54[4] = dm_int_st3_54[4];
	assign dm_int_st4_54[5] = dm_int_st3_54[5];
	assign dm_int_st4_54[6] = dm_int_st3_54[6];
	assign dm_int_st4_54[7] = dm_int_st3_54[7];
	assign dm_int_st4_54[8] = dm_int_st3_54[8];
	// Bit 55
	assign dm_int_st4_55[1] = dm_int_st3_55[0];
	assign dm_int_st4_55[2] = dm_int_st3_55[1];
	assign dm_int_st4_55[3] = dm_int_st3_55[2];
	assign dm_int_st4_55[4] = dm_int_st3_55[3];
	assign dm_int_st4_55[5] = dm_int_st3_55[4];
	assign dm_int_st4_55[6] = dm_int_st3_55[5];
	assign dm_int_st4_55[7] = dm_int_st3_55[6];
	assign dm_int_st4_55[8] = dm_int_st3_55[7];
	// Bit 56
	assign dm_int_st4_56[0] = dm_int_st3_56[0];
	assign dm_int_st4_56[1] = dm_int_st3_56[1];
	assign dm_int_st4_56[2] = dm_int_st3_56[2];
	assign dm_int_st4_56[3] = dm_int_st3_56[3];
	assign dm_int_st4_56[4] = dm_int_st3_56[4];
	assign dm_int_st4_56[5] = dm_int_st3_56[5];
	assign dm_int_st4_56[6] = dm_int_st3_56[6];
	// Bit 57
	assign dm_int_st4_57[0] = dm_int_st3_57[0];
	assign dm_int_st4_57[1] = dm_int_st3_57[1];
	assign dm_int_st4_57[2] = dm_int_st3_57[2];
	assign dm_int_st4_57[3] = dm_int_st3_57[3];
	assign dm_int_st4_57[4] = dm_int_st3_57[4];
	assign dm_int_st4_57[5] = dm_int_st3_57[5];
	// Bit 58
	assign dm_int_st4_58[0] = dm_int_st3_58[0];
	assign dm_int_st4_58[1] = dm_int_st3_58[1];
	assign dm_int_st4_58[2] = dm_int_st3_58[2];
	assign dm_int_st4_58[3] = dm_int_st3_58[3];
	assign dm_int_st4_58[4] = dm_int_st3_58[4];
	// Bit 59
	assign dm_int_st4_59[0] = dm_int_st3_59[0];
	assign dm_int_st4_59[1] = dm_int_st3_59[1];
	assign dm_int_st4_59[2] = dm_int_st3_59[2];
	assign dm_int_st4_59[3] = dm_int_st3_59[3];
	// Bit 60
	assign dm_int_st4_60[0] = dm_int_st3_60[0];
	assign dm_int_st4_60[1] = dm_int_st3_60[1];
	assign dm_int_st4_60[2] = dm_int_st3_60[2];
	// Bit 61
	assign dm_int_st4_61[0] = dm_int_st3_61[0];
	assign dm_int_st4_61[1] = dm_int_st3_61[1];
	// Bit 62
	assign dm_int_st4_62[0] = dm_int_st3_62[0];

	//// Stage 5 ////
	wire [0:0] dm_int_st5_0;
	wire [1:0] dm_int_st5_1;
	wire [2:0] dm_int_st5_2;
	wire [3:0] dm_int_st5_3;
	wire [4:0] dm_int_st5_4;
	wire [5:0] dm_int_st5_5;
	wire [5:0] dm_int_st5_6;
	wire [5:0] dm_int_st5_7;
	wire [5:0] dm_int_st5_8;
	wire [5:0] dm_int_st5_9;
	wire [5:0] dm_int_st5_10;
	wire [5:0] dm_int_st5_11;
	wire [5:0] dm_int_st5_12;
	wire [5:0] dm_int_st5_13;
	wire [5:0] dm_int_st5_14;
	wire [5:0] dm_int_st5_15;
	wire [5:0] dm_int_st5_16;
	wire [5:0] dm_int_st5_17;
	wire [5:0] dm_int_st5_18;
	wire [5:0] dm_int_st5_19;
	wire [5:0] dm_int_st5_20;
	wire [5:0] dm_int_st5_21;
	wire [5:0] dm_int_st5_22;
	wire [5:0] dm_int_st5_23;
	wire [5:0] dm_int_st5_24;
	wire [5:0] dm_int_st5_25;
	wire [5:0] dm_int_st5_26;
	wire [5:0] dm_int_st5_27;
	wire [5:0] dm_int_st5_28;
	wire [5:0] dm_int_st5_29;
	wire [5:0] dm_int_st5_30;
	wire [5:0] dm_int_st5_31;
	wire [5:0] dm_int_st5_32;
	wire [5:0] dm_int_st5_33;
	wire [5:0] dm_int_st5_34;
	wire [5:0] dm_int_st5_35;
	wire [5:0] dm_int_st5_36;
	wire [5:0] dm_int_st5_37;
	wire [5:0] dm_int_st5_38;
	wire [5:0] dm_int_st5_39;
	wire [5:0] dm_int_st5_40;
	wire [5:0] dm_int_st5_41;
	wire [5:0] dm_int_st5_42;
	wire [5:0] dm_int_st5_43;
	wire [5:0] dm_int_st5_44;
	wire [5:0] dm_int_st5_45;
	wire [5:0] dm_int_st5_46;
	wire [5:0] dm_int_st5_47;
	wire [5:0] dm_int_st5_48;
	wire [5:0] dm_int_st5_49;
	wire [5:0] dm_int_st5_50;
	wire [5:0] dm_int_st5_51;
	wire [5:0] dm_int_st5_52;
	wire [5:0] dm_int_st5_53;
	wire [5:0] dm_int_st5_54;
	wire [5:0] dm_int_st5_55;
	wire [5:0] dm_int_st5_56;
	wire [5:0] dm_int_st5_57;
	wire [5:0] dm_int_st5_58;
	wire [3:0] dm_int_st5_59;
	wire [2:0] dm_int_st5_60;
	wire [1:0] dm_int_st5_61;
	wire [0:0] dm_int_st5_62;

	// Bit 0
	assign dm_int_st5_0[0] = dm_int_st4_0[0];
	// Bit 1
	assign dm_int_st5_1[0] = dm_int_st4_1[0];
	assign dm_int_st5_1[1] = dm_int_st4_1[1];
	// Bit 2
	assign dm_int_st5_2[0] = dm_int_st4_2[0];
	assign dm_int_st5_2[1] = dm_int_st4_2[1];
	assign dm_int_st5_2[2] = dm_int_st4_2[2];
	// Bit 3
	assign dm_int_st5_3[0] = dm_int_st4_3[0];
	assign dm_int_st5_3[1] = dm_int_st4_3[1];
	assign dm_int_st5_3[2] = dm_int_st4_3[2];
	assign dm_int_st5_3[3] = dm_int_st4_3[3];
	// Bit 4
	assign dm_int_st5_4[0] = dm_int_st4_4[0];
	assign dm_int_st5_4[1] = dm_int_st4_4[1];
	assign dm_int_st5_4[2] = dm_int_st4_4[2];
	assign dm_int_st5_4[3] = dm_int_st4_4[3];
	assign dm_int_st5_4[4] = dm_int_st4_4[4];
	// Bit 5
	assign dm_int_st5_5[0] = dm_int_st4_5[0];
	assign dm_int_st5_5[1] = dm_int_st4_5[1];
	assign dm_int_st5_5[2] = dm_int_st4_5[2];
	assign dm_int_st5_5[3] = dm_int_st4_5[3];
	assign dm_int_st5_5[4] = dm_int_st4_5[4];
	assign dm_int_st5_5[5] = dm_int_st4_5[5];
	// Bit 6
	half_adder HA24(.a(dm_int_st4_6[0]), .b(dm_int_st4_6[1]), .s(dm_int_st5_6[0]), .cout(dm_int_st5_7[0]));
	assign dm_int_st5_6[1] = dm_int_st4_6[2];
	assign dm_int_st5_6[2] = dm_int_st4_6[3];
	assign dm_int_st5_6[3] = dm_int_st4_6[4];
	assign dm_int_st5_6[4] = dm_int_st4_6[5];
	assign dm_int_st5_6[5] = dm_int_st4_6[6];
	// Bit 7
	full_adder FA528(.a(dm_int_st4_7[0]), .b(dm_int_st4_7[1]), .cin(dm_int_st4_7[2]), .s(dm_int_st5_7[1]), .cout(dm_int_st5_8[0]));
	half_adder HA25(.a(dm_int_st4_7[3]), .b(dm_int_st4_7[4]), .s(dm_int_st5_7[2]), .cout(dm_int_st5_8[1]));
	assign dm_int_st5_7[3] = dm_int_st4_7[5];
	assign dm_int_st5_7[4] = dm_int_st4_7[6];
	assign dm_int_st5_7[5] = dm_int_st4_7[7];
	// Bit 8
	full_adder FA529(.a(dm_int_st4_8[0]), .b(dm_int_st4_8[1]), .cin(dm_int_st4_8[2]), .s(dm_int_st5_8[2]), .cout(dm_int_st5_9[0]));
	full_adder FA530(.a(dm_int_st4_8[3]), .b(dm_int_st4_8[4]), .cin(dm_int_st4_8[5]), .s(dm_int_st5_8[3]), .cout(dm_int_st5_9[1]));
	half_adder HA26(.a(dm_int_st4_8[6]), .b(dm_int_st4_8[7]), .s(dm_int_st5_8[4]), .cout(dm_int_st5_9[2]));
	assign dm_int_st5_8[5] = dm_int_st4_8[8];
	// Bit 9
	full_adder FA531(.a(dm_int_st4_9[0]), .b(dm_int_st4_9[1]), .cin(dm_int_st4_9[2]), .s(dm_int_st5_9[3]), .cout(dm_int_st5_10[0]));
	full_adder FA532(.a(dm_int_st4_9[3]), .b(dm_int_st4_9[4]), .cin(dm_int_st4_9[5]), .s(dm_int_st5_9[4]), .cout(dm_int_st5_10[1]));
	full_adder FA533(.a(dm_int_st4_9[6]), .b(dm_int_st4_9[7]), .cin(dm_int_st4_9[8]), .s(dm_int_st5_9[5]), .cout(dm_int_st5_10[2]));
	// Bit 10
	full_adder FA534(.a(dm_int_st4_10[0]), .b(dm_int_st4_10[1]), .cin(dm_int_st4_10[2]), .s(dm_int_st5_10[3]), .cout(dm_int_st5_11[0]));
	full_adder FA535(.a(dm_int_st4_10[3]), .b(dm_int_st4_10[4]), .cin(dm_int_st4_10[5]), .s(dm_int_st5_10[4]), .cout(dm_int_st5_11[1]));
	full_adder FA536(.a(dm_int_st4_10[6]), .b(dm_int_st4_10[7]), .cin(dm_int_st4_10[8]), .s(dm_int_st5_10[5]), .cout(dm_int_st5_11[2]));
	// Bit 11
	full_adder FA537(.a(dm_int_st4_11[0]), .b(dm_int_st4_11[1]), .cin(dm_int_st4_11[2]), .s(dm_int_st5_11[3]), .cout(dm_int_st5_12[0]));
	full_adder FA538(.a(dm_int_st4_11[3]), .b(dm_int_st4_11[4]), .cin(dm_int_st4_11[5]), .s(dm_int_st5_11[4]), .cout(dm_int_st5_12[1]));
	full_adder FA539(.a(dm_int_st4_11[6]), .b(dm_int_st4_11[7]), .cin(dm_int_st4_11[8]), .s(dm_int_st5_11[5]), .cout(dm_int_st5_12[2]));
	// Bit 12
	full_adder FA540(.a(dm_int_st4_12[0]), .b(dm_int_st4_12[1]), .cin(dm_int_st4_12[2]), .s(dm_int_st5_12[3]), .cout(dm_int_st5_13[0]));
	full_adder FA541(.a(dm_int_st4_12[3]), .b(dm_int_st4_12[4]), .cin(dm_int_st4_12[5]), .s(dm_int_st5_12[4]), .cout(dm_int_st5_13[1]));
	full_adder FA542(.a(dm_int_st4_12[6]), .b(dm_int_st4_12[7]), .cin(dm_int_st4_12[8]), .s(dm_int_st5_12[5]), .cout(dm_int_st5_13[2]));
	// Bit 13
	full_adder FA543(.a(dm_int_st4_13[0]), .b(dm_int_st4_13[1]), .cin(dm_int_st4_13[2]), .s(dm_int_st5_13[3]), .cout(dm_int_st5_14[0]));
	full_adder FA544(.a(dm_int_st4_13[3]), .b(dm_int_st4_13[4]), .cin(dm_int_st4_13[5]), .s(dm_int_st5_13[4]), .cout(dm_int_st5_14[1]));
	full_adder FA545(.a(dm_int_st4_13[6]), .b(dm_int_st4_13[7]), .cin(dm_int_st4_13[8]), .s(dm_int_st5_13[5]), .cout(dm_int_st5_14[2]));
	// Bit 14
	full_adder FA546(.a(dm_int_st4_14[0]), .b(dm_int_st4_14[1]), .cin(dm_int_st4_14[2]), .s(dm_int_st5_14[3]), .cout(dm_int_st5_15[0]));
	full_adder FA547(.a(dm_int_st4_14[3]), .b(dm_int_st4_14[4]), .cin(dm_int_st4_14[5]), .s(dm_int_st5_14[4]), .cout(dm_int_st5_15[1]));
	full_adder FA548(.a(dm_int_st4_14[6]), .b(dm_int_st4_14[7]), .cin(dm_int_st4_14[8]), .s(dm_int_st5_14[5]), .cout(dm_int_st5_15[2]));
	// Bit 15
	full_adder FA549(.a(dm_int_st4_15[0]), .b(dm_int_st4_15[1]), .cin(dm_int_st4_15[2]), .s(dm_int_st5_15[3]), .cout(dm_int_st5_16[0]));
	full_adder FA550(.a(dm_int_st4_15[3]), .b(dm_int_st4_15[4]), .cin(dm_int_st4_15[5]), .s(dm_int_st5_15[4]), .cout(dm_int_st5_16[1]));
	full_adder FA551(.a(dm_int_st4_15[6]), .b(dm_int_st4_15[7]), .cin(dm_int_st4_15[8]), .s(dm_int_st5_15[5]), .cout(dm_int_st5_16[2]));
	// Bit 16
	full_adder FA552(.a(dm_int_st4_16[0]), .b(dm_int_st4_16[1]), .cin(dm_int_st4_16[2]), .s(dm_int_st5_16[3]), .cout(dm_int_st5_17[0]));
	full_adder FA553(.a(dm_int_st4_16[3]), .b(dm_int_st4_16[4]), .cin(dm_int_st4_16[5]), .s(dm_int_st5_16[4]), .cout(dm_int_st5_17[1]));
	full_adder FA554(.a(dm_int_st4_16[6]), .b(dm_int_st4_16[7]), .cin(dm_int_st4_16[8]), .s(dm_int_st5_16[5]), .cout(dm_int_st5_17[2]));
	// Bit 17
	full_adder FA555(.a(dm_int_st4_17[0]), .b(dm_int_st4_17[1]), .cin(dm_int_st4_17[2]), .s(dm_int_st5_17[3]), .cout(dm_int_st5_18[0]));
	full_adder FA556(.a(dm_int_st4_17[3]), .b(dm_int_st4_17[4]), .cin(dm_int_st4_17[5]), .s(dm_int_st5_17[4]), .cout(dm_int_st5_18[1]));
	full_adder FA557(.a(dm_int_st4_17[6]), .b(dm_int_st4_17[7]), .cin(dm_int_st4_17[8]), .s(dm_int_st5_17[5]), .cout(dm_int_st5_18[2]));
	// Bit 18
	full_adder FA558(.a(dm_int_st4_18[0]), .b(dm_int_st4_18[1]), .cin(dm_int_st4_18[2]), .s(dm_int_st5_18[3]), .cout(dm_int_st5_19[0]));
	full_adder FA559(.a(dm_int_st4_18[3]), .b(dm_int_st4_18[4]), .cin(dm_int_st4_18[5]), .s(dm_int_st5_18[4]), .cout(dm_int_st5_19[1]));
	full_adder FA560(.a(dm_int_st4_18[6]), .b(dm_int_st4_18[7]), .cin(dm_int_st4_18[8]), .s(dm_int_st5_18[5]), .cout(dm_int_st5_19[2]));
	// Bit 19
	full_adder FA561(.a(dm_int_st4_19[0]), .b(dm_int_st4_19[1]), .cin(dm_int_st4_19[2]), .s(dm_int_st5_19[3]), .cout(dm_int_st5_20[0]));
	full_adder FA562(.a(dm_int_st4_19[3]), .b(dm_int_st4_19[4]), .cin(dm_int_st4_19[5]), .s(dm_int_st5_19[4]), .cout(dm_int_st5_20[1]));
	full_adder FA563(.a(dm_int_st4_19[6]), .b(dm_int_st4_19[7]), .cin(dm_int_st4_19[8]), .s(dm_int_st5_19[5]), .cout(dm_int_st5_20[2]));
	// Bit 20
	full_adder FA564(.a(dm_int_st4_20[0]), .b(dm_int_st4_20[1]), .cin(dm_int_st4_20[2]), .s(dm_int_st5_20[3]), .cout(dm_int_st5_21[0]));
	full_adder FA565(.a(dm_int_st4_20[3]), .b(dm_int_st4_20[4]), .cin(dm_int_st4_20[5]), .s(dm_int_st5_20[4]), .cout(dm_int_st5_21[1]));
	full_adder FA566(.a(dm_int_st4_20[6]), .b(dm_int_st4_20[7]), .cin(dm_int_st4_20[8]), .s(dm_int_st5_20[5]), .cout(dm_int_st5_21[2]));
	// Bit 21
	full_adder FA567(.a(dm_int_st4_21[0]), .b(dm_int_st4_21[1]), .cin(dm_int_st4_21[2]), .s(dm_int_st5_21[3]), .cout(dm_int_st5_22[0]));
	full_adder FA568(.a(dm_int_st4_21[3]), .b(dm_int_st4_21[4]), .cin(dm_int_st4_21[5]), .s(dm_int_st5_21[4]), .cout(dm_int_st5_22[1]));
	full_adder FA569(.a(dm_int_st4_21[6]), .b(dm_int_st4_21[7]), .cin(dm_int_st4_21[8]), .s(dm_int_st5_21[5]), .cout(dm_int_st5_22[2]));
	// Bit 22
	full_adder FA570(.a(dm_int_st4_22[0]), .b(dm_int_st4_22[1]), .cin(dm_int_st4_22[2]), .s(dm_int_st5_22[3]), .cout(dm_int_st5_23[0]));
	full_adder FA571(.a(dm_int_st4_22[3]), .b(dm_int_st4_22[4]), .cin(dm_int_st4_22[5]), .s(dm_int_st5_22[4]), .cout(dm_int_st5_23[1]));
	full_adder FA572(.a(dm_int_st4_22[6]), .b(dm_int_st4_22[7]), .cin(dm_int_st4_22[8]), .s(dm_int_st5_22[5]), .cout(dm_int_st5_23[2]));
	// Bit 23
	full_adder FA573(.a(dm_int_st4_23[0]), .b(dm_int_st4_23[1]), .cin(dm_int_st4_23[2]), .s(dm_int_st5_23[3]), .cout(dm_int_st5_24[0]));
	full_adder FA574(.a(dm_int_st4_23[3]), .b(dm_int_st4_23[4]), .cin(dm_int_st4_23[5]), .s(dm_int_st5_23[4]), .cout(dm_int_st5_24[1]));
	full_adder FA575(.a(dm_int_st4_23[6]), .b(dm_int_st4_23[7]), .cin(dm_int_st4_23[8]), .s(dm_int_st5_23[5]), .cout(dm_int_st5_24[2]));
	// Bit 24
	full_adder FA576(.a(dm_int_st4_24[0]), .b(dm_int_st4_24[1]), .cin(dm_int_st4_24[2]), .s(dm_int_st5_24[3]), .cout(dm_int_st5_25[0]));
	full_adder FA577(.a(dm_int_st4_24[3]), .b(dm_int_st4_24[4]), .cin(dm_int_st4_24[5]), .s(dm_int_st5_24[4]), .cout(dm_int_st5_25[1]));
	full_adder FA578(.a(dm_int_st4_24[6]), .b(dm_int_st4_24[7]), .cin(dm_int_st4_24[8]), .s(dm_int_st5_24[5]), .cout(dm_int_st5_25[2]));
	// Bit 25
	full_adder FA579(.a(dm_int_st4_25[0]), .b(dm_int_st4_25[1]), .cin(dm_int_st4_25[2]), .s(dm_int_st5_25[3]), .cout(dm_int_st5_26[0]));
	full_adder FA580(.a(dm_int_st4_25[3]), .b(dm_int_st4_25[4]), .cin(dm_int_st4_25[5]), .s(dm_int_st5_25[4]), .cout(dm_int_st5_26[1]));
	full_adder FA581(.a(dm_int_st4_25[6]), .b(dm_int_st4_25[7]), .cin(dm_int_st4_25[8]), .s(dm_int_st5_25[5]), .cout(dm_int_st5_26[2]));
	// Bit 26
	full_adder FA582(.a(dm_int_st4_26[0]), .b(dm_int_st4_26[1]), .cin(dm_int_st4_26[2]), .s(dm_int_st5_26[3]), .cout(dm_int_st5_27[0]));
	full_adder FA583(.a(dm_int_st4_26[3]), .b(dm_int_st4_26[4]), .cin(dm_int_st4_26[5]), .s(dm_int_st5_26[4]), .cout(dm_int_st5_27[1]));
	full_adder FA584(.a(dm_int_st4_26[6]), .b(dm_int_st4_26[7]), .cin(dm_int_st4_26[8]), .s(dm_int_st5_26[5]), .cout(dm_int_st5_27[2]));
	// Bit 27
	full_adder FA585(.a(dm_int_st4_27[0]), .b(dm_int_st4_27[1]), .cin(dm_int_st4_27[2]), .s(dm_int_st5_27[3]), .cout(dm_int_st5_28[0]));
	full_adder FA586(.a(dm_int_st4_27[3]), .b(dm_int_st4_27[4]), .cin(dm_int_st4_27[5]), .s(dm_int_st5_27[4]), .cout(dm_int_st5_28[1]));
	full_adder FA587(.a(dm_int_st4_27[6]), .b(dm_int_st4_27[7]), .cin(dm_int_st4_27[8]), .s(dm_int_st5_27[5]), .cout(dm_int_st5_28[2]));
	// Bit 28
	full_adder FA588(.a(dm_int_st4_28[0]), .b(dm_int_st4_28[1]), .cin(dm_int_st4_28[2]), .s(dm_int_st5_28[3]), .cout(dm_int_st5_29[0]));
	full_adder FA589(.a(dm_int_st4_28[3]), .b(dm_int_st4_28[4]), .cin(dm_int_st4_28[5]), .s(dm_int_st5_28[4]), .cout(dm_int_st5_29[1]));
	full_adder FA590(.a(dm_int_st4_28[6]), .b(dm_int_st4_28[7]), .cin(dm_int_st4_28[8]), .s(dm_int_st5_28[5]), .cout(dm_int_st5_29[2]));
	// Bit 29
	full_adder FA591(.a(dm_int_st4_29[0]), .b(dm_int_st4_29[1]), .cin(dm_int_st4_29[2]), .s(dm_int_st5_29[3]), .cout(dm_int_st5_30[0]));
	full_adder FA592(.a(dm_int_st4_29[3]), .b(dm_int_st4_29[4]), .cin(dm_int_st4_29[5]), .s(dm_int_st5_29[4]), .cout(dm_int_st5_30[1]));
	full_adder FA593(.a(dm_int_st4_29[6]), .b(dm_int_st4_29[7]), .cin(dm_int_st4_29[8]), .s(dm_int_st5_29[5]), .cout(dm_int_st5_30[2]));
	// Bit 30
	full_adder FA594(.a(dm_int_st4_30[0]), .b(dm_int_st4_30[1]), .cin(dm_int_st4_30[2]), .s(dm_int_st5_30[3]), .cout(dm_int_st5_31[0]));
	full_adder FA595(.a(dm_int_st4_30[3]), .b(dm_int_st4_30[4]), .cin(dm_int_st4_30[5]), .s(dm_int_st5_30[4]), .cout(dm_int_st5_31[1]));
	full_adder FA596(.a(dm_int_st4_30[6]), .b(dm_int_st4_30[7]), .cin(dm_int_st4_30[8]), .s(dm_int_st5_30[5]), .cout(dm_int_st5_31[2]));
	// Bit 31
	full_adder FA597(.a(dm_int_st4_31[0]), .b(dm_int_st4_31[1]), .cin(dm_int_st4_31[2]), .s(dm_int_st5_31[3]), .cout(dm_int_st5_32[0]));
	full_adder FA598(.a(dm_int_st4_31[3]), .b(dm_int_st4_31[4]), .cin(dm_int_st4_31[5]), .s(dm_int_st5_31[4]), .cout(dm_int_st5_32[1]));
	full_adder FA599(.a(dm_int_st4_31[6]), .b(dm_int_st4_31[7]), .cin(dm_int_st4_31[8]), .s(dm_int_st5_31[5]), .cout(dm_int_st5_32[2]));
	// Bit 32
	full_adder FA600(.a(dm_int_st4_32[0]), .b(dm_int_st4_32[1]), .cin(dm_int_st4_32[2]), .s(dm_int_st5_32[3]), .cout(dm_int_st5_33[0]));
	full_adder FA601(.a(dm_int_st4_32[3]), .b(dm_int_st4_32[4]), .cin(dm_int_st4_32[5]), .s(dm_int_st5_32[4]), .cout(dm_int_st5_33[1]));
	full_adder FA602(.a(dm_int_st4_32[6]), .b(dm_int_st4_32[7]), .cin(dm_int_st4_32[8]), .s(dm_int_st5_32[5]), .cout(dm_int_st5_33[2]));
	// Bit 33
	full_adder FA603(.a(dm_int_st4_33[0]), .b(dm_int_st4_33[1]), .cin(dm_int_st4_33[2]), .s(dm_int_st5_33[3]), .cout(dm_int_st5_34[0]));
	full_adder FA604(.a(dm_int_st4_33[3]), .b(dm_int_st4_33[4]), .cin(dm_int_st4_33[5]), .s(dm_int_st5_33[4]), .cout(dm_int_st5_34[1]));
	full_adder FA605(.a(dm_int_st4_33[6]), .b(dm_int_st4_33[7]), .cin(dm_int_st4_33[8]), .s(dm_int_st5_33[5]), .cout(dm_int_st5_34[2]));
	// Bit 34
	full_adder FA606(.a(dm_int_st4_34[0]), .b(dm_int_st4_34[1]), .cin(dm_int_st4_34[2]), .s(dm_int_st5_34[3]), .cout(dm_int_st5_35[0]));
	full_adder FA607(.a(dm_int_st4_34[3]), .b(dm_int_st4_34[4]), .cin(dm_int_st4_34[5]), .s(dm_int_st5_34[4]), .cout(dm_int_st5_35[1]));
	full_adder FA608(.a(dm_int_st4_34[6]), .b(dm_int_st4_34[7]), .cin(dm_int_st4_34[8]), .s(dm_int_st5_34[5]), .cout(dm_int_st5_35[2]));
	// Bit 35
	full_adder FA609(.a(dm_int_st4_35[0]), .b(dm_int_st4_35[1]), .cin(dm_int_st4_35[2]), .s(dm_int_st5_35[3]), .cout(dm_int_st5_36[0]));
	full_adder FA610(.a(dm_int_st4_35[3]), .b(dm_int_st4_35[4]), .cin(dm_int_st4_35[5]), .s(dm_int_st5_35[4]), .cout(dm_int_st5_36[1]));
	full_adder FA611(.a(dm_int_st4_35[6]), .b(dm_int_st4_35[7]), .cin(dm_int_st4_35[8]), .s(dm_int_st5_35[5]), .cout(dm_int_st5_36[2]));
	// Bit 36
	full_adder FA612(.a(dm_int_st4_36[0]), .b(dm_int_st4_36[1]), .cin(dm_int_st4_36[2]), .s(dm_int_st5_36[3]), .cout(dm_int_st5_37[0]));
	full_adder FA613(.a(dm_int_st4_36[3]), .b(dm_int_st4_36[4]), .cin(dm_int_st4_36[5]), .s(dm_int_st5_36[4]), .cout(dm_int_st5_37[1]));
	full_adder FA614(.a(dm_int_st4_36[6]), .b(dm_int_st4_36[7]), .cin(dm_int_st4_36[8]), .s(dm_int_st5_36[5]), .cout(dm_int_st5_37[2]));
	// Bit 37
	full_adder FA615(.a(dm_int_st4_37[0]), .b(dm_int_st4_37[1]), .cin(dm_int_st4_37[2]), .s(dm_int_st5_37[3]), .cout(dm_int_st5_38[0]));
	full_adder FA616(.a(dm_int_st4_37[3]), .b(dm_int_st4_37[4]), .cin(dm_int_st4_37[5]), .s(dm_int_st5_37[4]), .cout(dm_int_st5_38[1]));
	full_adder FA617(.a(dm_int_st4_37[6]), .b(dm_int_st4_37[7]), .cin(dm_int_st4_37[8]), .s(dm_int_st5_37[5]), .cout(dm_int_st5_38[2]));
	// Bit 38
	full_adder FA618(.a(dm_int_st4_38[0]), .b(dm_int_st4_38[1]), .cin(dm_int_st4_38[2]), .s(dm_int_st5_38[3]), .cout(dm_int_st5_39[0]));
	full_adder FA619(.a(dm_int_st4_38[3]), .b(dm_int_st4_38[4]), .cin(dm_int_st4_38[5]), .s(dm_int_st5_38[4]), .cout(dm_int_st5_39[1]));
	full_adder FA620(.a(dm_int_st4_38[6]), .b(dm_int_st4_38[7]), .cin(dm_int_st4_38[8]), .s(dm_int_st5_38[5]), .cout(dm_int_st5_39[2]));
	// Bit 39
	full_adder FA621(.a(dm_int_st4_39[0]), .b(dm_int_st4_39[1]), .cin(dm_int_st4_39[2]), .s(dm_int_st5_39[3]), .cout(dm_int_st5_40[0]));
	full_adder FA622(.a(dm_int_st4_39[3]), .b(dm_int_st4_39[4]), .cin(dm_int_st4_39[5]), .s(dm_int_st5_39[4]), .cout(dm_int_st5_40[1]));
	full_adder FA623(.a(dm_int_st4_39[6]), .b(dm_int_st4_39[7]), .cin(dm_int_st4_39[8]), .s(dm_int_st5_39[5]), .cout(dm_int_st5_40[2]));
	// Bit 40
	full_adder FA624(.a(dm_int_st4_40[0]), .b(dm_int_st4_40[1]), .cin(dm_int_st4_40[2]), .s(dm_int_st5_40[3]), .cout(dm_int_st5_41[0]));
	full_adder FA625(.a(dm_int_st4_40[3]), .b(dm_int_st4_40[4]), .cin(dm_int_st4_40[5]), .s(dm_int_st5_40[4]), .cout(dm_int_st5_41[1]));
	full_adder FA626(.a(dm_int_st4_40[6]), .b(dm_int_st4_40[7]), .cin(dm_int_st4_40[8]), .s(dm_int_st5_40[5]), .cout(dm_int_st5_41[2]));
	// Bit 41
	full_adder FA627(.a(dm_int_st4_41[0]), .b(dm_int_st4_41[1]), .cin(dm_int_st4_41[2]), .s(dm_int_st5_41[3]), .cout(dm_int_st5_42[0]));
	full_adder FA628(.a(dm_int_st4_41[3]), .b(dm_int_st4_41[4]), .cin(dm_int_st4_41[5]), .s(dm_int_st5_41[4]), .cout(dm_int_st5_42[1]));
	full_adder FA629(.a(dm_int_st4_41[6]), .b(dm_int_st4_41[7]), .cin(dm_int_st4_41[8]), .s(dm_int_st5_41[5]), .cout(dm_int_st5_42[2]));
	// Bit 42
	full_adder FA630(.a(dm_int_st4_42[0]), .b(dm_int_st4_42[1]), .cin(dm_int_st4_42[2]), .s(dm_int_st5_42[3]), .cout(dm_int_st5_43[0]));
	full_adder FA631(.a(dm_int_st4_42[3]), .b(dm_int_st4_42[4]), .cin(dm_int_st4_42[5]), .s(dm_int_st5_42[4]), .cout(dm_int_st5_43[1]));
	full_adder FA632(.a(dm_int_st4_42[6]), .b(dm_int_st4_42[7]), .cin(dm_int_st4_42[8]), .s(dm_int_st5_42[5]), .cout(dm_int_st5_43[2]));
	// Bit 43
	full_adder FA633(.a(dm_int_st4_43[0]), .b(dm_int_st4_43[1]), .cin(dm_int_st4_43[2]), .s(dm_int_st5_43[3]), .cout(dm_int_st5_44[0]));
	full_adder FA634(.a(dm_int_st4_43[3]), .b(dm_int_st4_43[4]), .cin(dm_int_st4_43[5]), .s(dm_int_st5_43[4]), .cout(dm_int_st5_44[1]));
	full_adder FA635(.a(dm_int_st4_43[6]), .b(dm_int_st4_43[7]), .cin(dm_int_st4_43[8]), .s(dm_int_st5_43[5]), .cout(dm_int_st5_44[2]));
	// Bit 44
	full_adder FA636(.a(dm_int_st4_44[0]), .b(dm_int_st4_44[1]), .cin(dm_int_st4_44[2]), .s(dm_int_st5_44[3]), .cout(dm_int_st5_45[0]));
	full_adder FA637(.a(dm_int_st4_44[3]), .b(dm_int_st4_44[4]), .cin(dm_int_st4_44[5]), .s(dm_int_st5_44[4]), .cout(dm_int_st5_45[1]));
	full_adder FA638(.a(dm_int_st4_44[6]), .b(dm_int_st4_44[7]), .cin(dm_int_st4_44[8]), .s(dm_int_st5_44[5]), .cout(dm_int_st5_45[2]));
	// Bit 45
	full_adder FA639(.a(dm_int_st4_45[0]), .b(dm_int_st4_45[1]), .cin(dm_int_st4_45[2]), .s(dm_int_st5_45[3]), .cout(dm_int_st5_46[0]));
	full_adder FA640(.a(dm_int_st4_45[3]), .b(dm_int_st4_45[4]), .cin(dm_int_st4_45[5]), .s(dm_int_st5_45[4]), .cout(dm_int_st5_46[1]));
	full_adder FA641(.a(dm_int_st4_45[6]), .b(dm_int_st4_45[7]), .cin(dm_int_st4_45[8]), .s(dm_int_st5_45[5]), .cout(dm_int_st5_46[2]));
	// Bit 46
	full_adder FA642(.a(dm_int_st4_46[0]), .b(dm_int_st4_46[1]), .cin(dm_int_st4_46[2]), .s(dm_int_st5_46[3]), .cout(dm_int_st5_47[0]));
	full_adder FA643(.a(dm_int_st4_46[3]), .b(dm_int_st4_46[4]), .cin(dm_int_st4_46[5]), .s(dm_int_st5_46[4]), .cout(dm_int_st5_47[1]));
	full_adder FA644(.a(dm_int_st4_46[6]), .b(dm_int_st4_46[7]), .cin(dm_int_st4_46[8]), .s(dm_int_st5_46[5]), .cout(dm_int_st5_47[2]));
	// Bit 47
	full_adder FA645(.a(dm_int_st4_47[0]), .b(dm_int_st4_47[1]), .cin(dm_int_st4_47[2]), .s(dm_int_st5_47[3]), .cout(dm_int_st5_48[0]));
	full_adder FA646(.a(dm_int_st4_47[3]), .b(dm_int_st4_47[4]), .cin(dm_int_st4_47[5]), .s(dm_int_st5_47[4]), .cout(dm_int_st5_48[1]));
	full_adder FA647(.a(dm_int_st4_47[6]), .b(dm_int_st4_47[7]), .cin(dm_int_st4_47[8]), .s(dm_int_st5_47[5]), .cout(dm_int_st5_48[2]));
	// Bit 48
	full_adder FA648(.a(dm_int_st4_48[0]), .b(dm_int_st4_48[1]), .cin(dm_int_st4_48[2]), .s(dm_int_st5_48[3]), .cout(dm_int_st5_49[0]));
	full_adder FA649(.a(dm_int_st4_48[3]), .b(dm_int_st4_48[4]), .cin(dm_int_st4_48[5]), .s(dm_int_st5_48[4]), .cout(dm_int_st5_49[1]));
	full_adder FA650(.a(dm_int_st4_48[6]), .b(dm_int_st4_48[7]), .cin(dm_int_st4_48[8]), .s(dm_int_st5_48[5]), .cout(dm_int_st5_49[2]));
	// Bit 49
	full_adder FA651(.a(dm_int_st4_49[0]), .b(dm_int_st4_49[1]), .cin(dm_int_st4_49[2]), .s(dm_int_st5_49[3]), .cout(dm_int_st5_50[0]));
	full_adder FA652(.a(dm_int_st4_49[3]), .b(dm_int_st4_49[4]), .cin(dm_int_st4_49[5]), .s(dm_int_st5_49[4]), .cout(dm_int_st5_50[1]));
	full_adder FA653(.a(dm_int_st4_49[6]), .b(dm_int_st4_49[7]), .cin(dm_int_st4_49[8]), .s(dm_int_st5_49[5]), .cout(dm_int_st5_50[2]));
	// Bit 50
	full_adder FA654(.a(dm_int_st4_50[0]), .b(dm_int_st4_50[1]), .cin(dm_int_st4_50[2]), .s(dm_int_st5_50[3]), .cout(dm_int_st5_51[0]));
	full_adder FA655(.a(dm_int_st4_50[3]), .b(dm_int_st4_50[4]), .cin(dm_int_st4_50[5]), .s(dm_int_st5_50[4]), .cout(dm_int_st5_51[1]));
	full_adder FA656(.a(dm_int_st4_50[6]), .b(dm_int_st4_50[7]), .cin(dm_int_st4_50[8]), .s(dm_int_st5_50[5]), .cout(dm_int_st5_51[2]));
	// Bit 51
	full_adder FA657(.a(dm_int_st4_51[0]), .b(dm_int_st4_51[1]), .cin(dm_int_st4_51[2]), .s(dm_int_st5_51[3]), .cout(dm_int_st5_52[0]));
	full_adder FA658(.a(dm_int_st4_51[3]), .b(dm_int_st4_51[4]), .cin(dm_int_st4_51[5]), .s(dm_int_st5_51[4]), .cout(dm_int_st5_52[1]));
	full_adder FA659(.a(dm_int_st4_51[6]), .b(dm_int_st4_51[7]), .cin(dm_int_st4_51[8]), .s(dm_int_st5_51[5]), .cout(dm_int_st5_52[2]));
	// Bit 52
	full_adder FA660(.a(dm_int_st4_52[0]), .b(dm_int_st4_52[1]), .cin(dm_int_st4_52[2]), .s(dm_int_st5_52[3]), .cout(dm_int_st5_53[0]));
	full_adder FA661(.a(dm_int_st4_52[3]), .b(dm_int_st4_52[4]), .cin(dm_int_st4_52[5]), .s(dm_int_st5_52[4]), .cout(dm_int_st5_53[1]));
	full_adder FA662(.a(dm_int_st4_52[6]), .b(dm_int_st4_52[7]), .cin(dm_int_st4_52[8]), .s(dm_int_st5_52[5]), .cout(dm_int_st5_53[2]));
	// Bit 53
	full_adder FA663(.a(dm_int_st4_53[0]), .b(dm_int_st4_53[1]), .cin(dm_int_st4_53[2]), .s(dm_int_st5_53[3]), .cout(dm_int_st5_54[0]));
	full_adder FA664(.a(dm_int_st4_53[3]), .b(dm_int_st4_53[4]), .cin(dm_int_st4_53[5]), .s(dm_int_st5_53[4]), .cout(dm_int_st5_54[1]));
	full_adder FA665(.a(dm_int_st4_53[6]), .b(dm_int_st4_53[7]), .cin(dm_int_st4_53[8]), .s(dm_int_st5_53[5]), .cout(dm_int_st5_54[2]));
	// Bit 54
	full_adder FA666(.a(dm_int_st4_54[0]), .b(dm_int_st4_54[1]), .cin(dm_int_st4_54[2]), .s(dm_int_st5_54[3]), .cout(dm_int_st5_55[0]));
	full_adder FA667(.a(dm_int_st4_54[3]), .b(dm_int_st4_54[4]), .cin(dm_int_st4_54[5]), .s(dm_int_st5_54[4]), .cout(dm_int_st5_55[1]));
	full_adder FA668(.a(dm_int_st4_54[6]), .b(dm_int_st4_54[7]), .cin(dm_int_st4_54[8]), .s(dm_int_st5_54[5]), .cout(dm_int_st5_55[2]));
	// Bit 55
	full_adder FA669(.a(dm_int_st4_55[0]), .b(dm_int_st4_55[1]), .cin(dm_int_st4_55[2]), .s(dm_int_st5_55[3]), .cout(dm_int_st5_56[0]));
	full_adder FA670(.a(dm_int_st4_55[3]), .b(dm_int_st4_55[4]), .cin(dm_int_st4_55[5]), .s(dm_int_st5_55[4]), .cout(dm_int_st5_56[1]));
	full_adder FA671(.a(dm_int_st4_55[6]), .b(dm_int_st4_55[7]), .cin(dm_int_st4_55[8]), .s(dm_int_st5_55[5]), .cout(dm_int_st5_56[2]));
	// Bit 56
	full_adder FA672(.a(dm_int_st4_56[0]), .b(dm_int_st4_56[1]), .cin(dm_int_st4_56[2]), .s(dm_int_st5_56[3]), .cout(dm_int_st5_57[0]));
	full_adder FA673(.a(dm_int_st4_56[3]), .b(dm_int_st4_56[4]), .cin(dm_int_st4_56[5]), .s(dm_int_st5_56[4]), .cout(dm_int_st5_57[1]));
	assign dm_int_st5_56[5] = dm_int_st4_56[6];
	// Bit 57
	full_adder FA674(.a(dm_int_st4_57[0]), .b(dm_int_st4_57[1]), .cin(dm_int_st4_57[2]), .s(dm_int_st5_57[2]), .cout(dm_int_st5_58[0]));
	assign dm_int_st5_57[3] = dm_int_st4_57[3];
	assign dm_int_st5_57[4] = dm_int_st4_57[4];
	assign dm_int_st5_57[5] = dm_int_st4_57[5];
	// Bit 58
	assign dm_int_st5_58[1] = dm_int_st4_58[0];
	assign dm_int_st5_58[2] = dm_int_st4_58[1];
	assign dm_int_st5_58[3] = dm_int_st4_58[2];
	assign dm_int_st5_58[4] = dm_int_st4_58[3];
	assign dm_int_st5_58[5] = dm_int_st4_58[4];
	// Bit 59
	assign dm_int_st5_59[0] = dm_int_st4_59[0];
	assign dm_int_st5_59[1] = dm_int_st4_59[1];
	assign dm_int_st5_59[2] = dm_int_st4_59[2];
	assign dm_int_st5_59[3] = dm_int_st4_59[3];
	// Bit 60
	assign dm_int_st5_60[0] = dm_int_st4_60[0];
	assign dm_int_st5_60[1] = dm_int_st4_60[1];
	assign dm_int_st5_60[2] = dm_int_st4_60[2];
	// Bit 61
	assign dm_int_st5_61[0] = dm_int_st4_61[0];
	assign dm_int_st5_61[1] = dm_int_st4_61[1];
	// Bit 62
	assign dm_int_st5_62[0] = dm_int_st4_62[0];

	//// Stage 6 ////
	wire [0:0] dm_int_st6_0;
	wire [1:0] dm_int_st6_1;
	wire [2:0] dm_int_st6_2;
	wire [3:0] dm_int_st6_3;
	wire [3:0] dm_int_st6_4;
	wire [3:0] dm_int_st6_5;
	wire [3:0] dm_int_st6_6;
	wire [3:0] dm_int_st6_7;
	wire [3:0] dm_int_st6_8;
	wire [3:0] dm_int_st6_9;
	wire [3:0] dm_int_st6_10;
	wire [3:0] dm_int_st6_11;
	wire [3:0] dm_int_st6_12;
	wire [3:0] dm_int_st6_13;
	wire [3:0] dm_int_st6_14;
	wire [3:0] dm_int_st6_15;
	wire [3:0] dm_int_st6_16;
	wire [3:0] dm_int_st6_17;
	wire [3:0] dm_int_st6_18;
	wire [3:0] dm_int_st6_19;
	wire [3:0] dm_int_st6_20;
	wire [3:0] dm_int_st6_21;
	wire [3:0] dm_int_st6_22;
	wire [3:0] dm_int_st6_23;
	wire [3:0] dm_int_st6_24;
	wire [3:0] dm_int_st6_25;
	wire [3:0] dm_int_st6_26;
	wire [3:0] dm_int_st6_27;
	wire [3:0] dm_int_st6_28;
	wire [3:0] dm_int_st6_29;
	wire [3:0] dm_int_st6_30;
	wire [3:0] dm_int_st6_31;
	wire [3:0] dm_int_st6_32;
	wire [3:0] dm_int_st6_33;
	wire [3:0] dm_int_st6_34;
	wire [3:0] dm_int_st6_35;
	wire [3:0] dm_int_st6_36;
	wire [3:0] dm_int_st6_37;
	wire [3:0] dm_int_st6_38;
	wire [3:0] dm_int_st6_39;
	wire [3:0] dm_int_st6_40;
	wire [3:0] dm_int_st6_41;
	wire [3:0] dm_int_st6_42;
	wire [3:0] dm_int_st6_43;
	wire [3:0] dm_int_st6_44;
	wire [3:0] dm_int_st6_45;
	wire [3:0] dm_int_st6_46;
	wire [3:0] dm_int_st6_47;
	wire [3:0] dm_int_st6_48;
	wire [3:0] dm_int_st6_49;
	wire [3:0] dm_int_st6_50;
	wire [3:0] dm_int_st6_51;
	wire [3:0] dm_int_st6_52;
	wire [3:0] dm_int_st6_53;
	wire [3:0] dm_int_st6_54;
	wire [3:0] dm_int_st6_55;
	wire [3:0] dm_int_st6_56;
	wire [3:0] dm_int_st6_57;
	wire [3:0] dm_int_st6_58;
	wire [3:0] dm_int_st6_59;
	wire [3:0] dm_int_st6_60;
	wire [1:0] dm_int_st6_61;
	wire [0:0] dm_int_st6_62;

	// Bit 0
	assign dm_int_st6_0[0] = dm_int_st5_0[0];
	// Bit 1
	assign dm_int_st6_1[0] = dm_int_st5_1[0];
	assign dm_int_st6_1[1] = dm_int_st5_1[1];
	// Bit 2
	assign dm_int_st6_2[0] = dm_int_st5_2[0];
	assign dm_int_st6_2[1] = dm_int_st5_2[1];
	assign dm_int_st6_2[2] = dm_int_st5_2[2];
	// Bit 3
	assign dm_int_st6_3[0] = dm_int_st5_3[0];
	assign dm_int_st6_3[1] = dm_int_st5_3[1];
	assign dm_int_st6_3[2] = dm_int_st5_3[2];
	assign dm_int_st6_3[3] = dm_int_st5_3[3];
	// Bit 4
	half_adder HA27(.a(dm_int_st5_4[0]), .b(dm_int_st5_4[1]), .s(dm_int_st6_4[0]), .cout(dm_int_st6_5[0]));
	assign dm_int_st6_4[1] = dm_int_st5_4[2];
	assign dm_int_st6_4[2] = dm_int_st5_4[3];
	assign dm_int_st6_4[3] = dm_int_st5_4[4];
	// Bit 5
	full_adder FA675(.a(dm_int_st5_5[0]), .b(dm_int_st5_5[1]), .cin(dm_int_st5_5[2]), .s(dm_int_st6_5[1]), .cout(dm_int_st6_6[0]));
	half_adder HA28(.a(dm_int_st5_5[3]), .b(dm_int_st5_5[4]), .s(dm_int_st6_5[2]), .cout(dm_int_st6_6[1]));
	assign dm_int_st6_5[3] = dm_int_st5_5[5];
	// Bit 6
	full_adder FA676(.a(dm_int_st5_6[0]), .b(dm_int_st5_6[1]), .cin(dm_int_st5_6[2]), .s(dm_int_st6_6[2]), .cout(dm_int_st6_7[0]));
	full_adder FA677(.a(dm_int_st5_6[3]), .b(dm_int_st5_6[4]), .cin(dm_int_st5_6[5]), .s(dm_int_st6_6[3]), .cout(dm_int_st6_7[1]));
	// Bit 7
	full_adder FA678(.a(dm_int_st5_7[0]), .b(dm_int_st5_7[1]), .cin(dm_int_st5_7[2]), .s(dm_int_st6_7[2]), .cout(dm_int_st6_8[0]));
	full_adder FA679(.a(dm_int_st5_7[3]), .b(dm_int_st5_7[4]), .cin(dm_int_st5_7[5]), .s(dm_int_st6_7[3]), .cout(dm_int_st6_8[1]));
	// Bit 8
	full_adder FA680(.a(dm_int_st5_8[0]), .b(dm_int_st5_8[1]), .cin(dm_int_st5_8[2]), .s(dm_int_st6_8[2]), .cout(dm_int_st6_9[0]));
	full_adder FA681(.a(dm_int_st5_8[3]), .b(dm_int_st5_8[4]), .cin(dm_int_st5_8[5]), .s(dm_int_st6_8[3]), .cout(dm_int_st6_9[1]));
	// Bit 9
	full_adder FA682(.a(dm_int_st5_9[0]), .b(dm_int_st5_9[1]), .cin(dm_int_st5_9[2]), .s(dm_int_st6_9[2]), .cout(dm_int_st6_10[0]));
	full_adder FA683(.a(dm_int_st5_9[3]), .b(dm_int_st5_9[4]), .cin(dm_int_st5_9[5]), .s(dm_int_st6_9[3]), .cout(dm_int_st6_10[1]));
	// Bit 10
	full_adder FA684(.a(dm_int_st5_10[0]), .b(dm_int_st5_10[1]), .cin(dm_int_st5_10[2]), .s(dm_int_st6_10[2]), .cout(dm_int_st6_11[0]));
	full_adder FA685(.a(dm_int_st5_10[3]), .b(dm_int_st5_10[4]), .cin(dm_int_st5_10[5]), .s(dm_int_st6_10[3]), .cout(dm_int_st6_11[1]));
	// Bit 11
	full_adder FA686(.a(dm_int_st5_11[0]), .b(dm_int_st5_11[1]), .cin(dm_int_st5_11[2]), .s(dm_int_st6_11[2]), .cout(dm_int_st6_12[0]));
	full_adder FA687(.a(dm_int_st5_11[3]), .b(dm_int_st5_11[4]), .cin(dm_int_st5_11[5]), .s(dm_int_st6_11[3]), .cout(dm_int_st6_12[1]));
	// Bit 12
	full_adder FA688(.a(dm_int_st5_12[0]), .b(dm_int_st5_12[1]), .cin(dm_int_st5_12[2]), .s(dm_int_st6_12[2]), .cout(dm_int_st6_13[0]));
	full_adder FA689(.a(dm_int_st5_12[3]), .b(dm_int_st5_12[4]), .cin(dm_int_st5_12[5]), .s(dm_int_st6_12[3]), .cout(dm_int_st6_13[1]));
	// Bit 13
	full_adder FA690(.a(dm_int_st5_13[0]), .b(dm_int_st5_13[1]), .cin(dm_int_st5_13[2]), .s(dm_int_st6_13[2]), .cout(dm_int_st6_14[0]));
	full_adder FA691(.a(dm_int_st5_13[3]), .b(dm_int_st5_13[4]), .cin(dm_int_st5_13[5]), .s(dm_int_st6_13[3]), .cout(dm_int_st6_14[1]));
	// Bit 14
	full_adder FA692(.a(dm_int_st5_14[0]), .b(dm_int_st5_14[1]), .cin(dm_int_st5_14[2]), .s(dm_int_st6_14[2]), .cout(dm_int_st6_15[0]));
	full_adder FA693(.a(dm_int_st5_14[3]), .b(dm_int_st5_14[4]), .cin(dm_int_st5_14[5]), .s(dm_int_st6_14[3]), .cout(dm_int_st6_15[1]));
	// Bit 15
	full_adder FA694(.a(dm_int_st5_15[0]), .b(dm_int_st5_15[1]), .cin(dm_int_st5_15[2]), .s(dm_int_st6_15[2]), .cout(dm_int_st6_16[0]));
	full_adder FA695(.a(dm_int_st5_15[3]), .b(dm_int_st5_15[4]), .cin(dm_int_st5_15[5]), .s(dm_int_st6_15[3]), .cout(dm_int_st6_16[1]));
	// Bit 16
	full_adder FA696(.a(dm_int_st5_16[0]), .b(dm_int_st5_16[1]), .cin(dm_int_st5_16[2]), .s(dm_int_st6_16[2]), .cout(dm_int_st6_17[0]));
	full_adder FA697(.a(dm_int_st5_16[3]), .b(dm_int_st5_16[4]), .cin(dm_int_st5_16[5]), .s(dm_int_st6_16[3]), .cout(dm_int_st6_17[1]));
	// Bit 17
	full_adder FA698(.a(dm_int_st5_17[0]), .b(dm_int_st5_17[1]), .cin(dm_int_st5_17[2]), .s(dm_int_st6_17[2]), .cout(dm_int_st6_18[0]));
	full_adder FA699(.a(dm_int_st5_17[3]), .b(dm_int_st5_17[4]), .cin(dm_int_st5_17[5]), .s(dm_int_st6_17[3]), .cout(dm_int_st6_18[1]));
	// Bit 18
	full_adder FA700(.a(dm_int_st5_18[0]), .b(dm_int_st5_18[1]), .cin(dm_int_st5_18[2]), .s(dm_int_st6_18[2]), .cout(dm_int_st6_19[0]));
	full_adder FA701(.a(dm_int_st5_18[3]), .b(dm_int_st5_18[4]), .cin(dm_int_st5_18[5]), .s(dm_int_st6_18[3]), .cout(dm_int_st6_19[1]));
	// Bit 19
	full_adder FA702(.a(dm_int_st5_19[0]), .b(dm_int_st5_19[1]), .cin(dm_int_st5_19[2]), .s(dm_int_st6_19[2]), .cout(dm_int_st6_20[0]));
	full_adder FA703(.a(dm_int_st5_19[3]), .b(dm_int_st5_19[4]), .cin(dm_int_st5_19[5]), .s(dm_int_st6_19[3]), .cout(dm_int_st6_20[1]));
	// Bit 20
	full_adder FA704(.a(dm_int_st5_20[0]), .b(dm_int_st5_20[1]), .cin(dm_int_st5_20[2]), .s(dm_int_st6_20[2]), .cout(dm_int_st6_21[0]));
	full_adder FA705(.a(dm_int_st5_20[3]), .b(dm_int_st5_20[4]), .cin(dm_int_st5_20[5]), .s(dm_int_st6_20[3]), .cout(dm_int_st6_21[1]));
	// Bit 21
	full_adder FA706(.a(dm_int_st5_21[0]), .b(dm_int_st5_21[1]), .cin(dm_int_st5_21[2]), .s(dm_int_st6_21[2]), .cout(dm_int_st6_22[0]));
	full_adder FA707(.a(dm_int_st5_21[3]), .b(dm_int_st5_21[4]), .cin(dm_int_st5_21[5]), .s(dm_int_st6_21[3]), .cout(dm_int_st6_22[1]));
	// Bit 22
	full_adder FA708(.a(dm_int_st5_22[0]), .b(dm_int_st5_22[1]), .cin(dm_int_st5_22[2]), .s(dm_int_st6_22[2]), .cout(dm_int_st6_23[0]));
	full_adder FA709(.a(dm_int_st5_22[3]), .b(dm_int_st5_22[4]), .cin(dm_int_st5_22[5]), .s(dm_int_st6_22[3]), .cout(dm_int_st6_23[1]));
	// Bit 23
	full_adder FA710(.a(dm_int_st5_23[0]), .b(dm_int_st5_23[1]), .cin(dm_int_st5_23[2]), .s(dm_int_st6_23[2]), .cout(dm_int_st6_24[0]));
	full_adder FA711(.a(dm_int_st5_23[3]), .b(dm_int_st5_23[4]), .cin(dm_int_st5_23[5]), .s(dm_int_st6_23[3]), .cout(dm_int_st6_24[1]));
	// Bit 24
	full_adder FA712(.a(dm_int_st5_24[0]), .b(dm_int_st5_24[1]), .cin(dm_int_st5_24[2]), .s(dm_int_st6_24[2]), .cout(dm_int_st6_25[0]));
	full_adder FA713(.a(dm_int_st5_24[3]), .b(dm_int_st5_24[4]), .cin(dm_int_st5_24[5]), .s(dm_int_st6_24[3]), .cout(dm_int_st6_25[1]));
	// Bit 25
	full_adder FA714(.a(dm_int_st5_25[0]), .b(dm_int_st5_25[1]), .cin(dm_int_st5_25[2]), .s(dm_int_st6_25[2]), .cout(dm_int_st6_26[0]));
	full_adder FA715(.a(dm_int_st5_25[3]), .b(dm_int_st5_25[4]), .cin(dm_int_st5_25[5]), .s(dm_int_st6_25[3]), .cout(dm_int_st6_26[1]));
	// Bit 26
	full_adder FA716(.a(dm_int_st5_26[0]), .b(dm_int_st5_26[1]), .cin(dm_int_st5_26[2]), .s(dm_int_st6_26[2]), .cout(dm_int_st6_27[0]));
	full_adder FA717(.a(dm_int_st5_26[3]), .b(dm_int_st5_26[4]), .cin(dm_int_st5_26[5]), .s(dm_int_st6_26[3]), .cout(dm_int_st6_27[1]));
	// Bit 27
	full_adder FA718(.a(dm_int_st5_27[0]), .b(dm_int_st5_27[1]), .cin(dm_int_st5_27[2]), .s(dm_int_st6_27[2]), .cout(dm_int_st6_28[0]));
	full_adder FA719(.a(dm_int_st5_27[3]), .b(dm_int_st5_27[4]), .cin(dm_int_st5_27[5]), .s(dm_int_st6_27[3]), .cout(dm_int_st6_28[1]));
	// Bit 28
	full_adder FA720(.a(dm_int_st5_28[0]), .b(dm_int_st5_28[1]), .cin(dm_int_st5_28[2]), .s(dm_int_st6_28[2]), .cout(dm_int_st6_29[0]));
	full_adder FA721(.a(dm_int_st5_28[3]), .b(dm_int_st5_28[4]), .cin(dm_int_st5_28[5]), .s(dm_int_st6_28[3]), .cout(dm_int_st6_29[1]));
	// Bit 29
	full_adder FA722(.a(dm_int_st5_29[0]), .b(dm_int_st5_29[1]), .cin(dm_int_st5_29[2]), .s(dm_int_st6_29[2]), .cout(dm_int_st6_30[0]));
	full_adder FA723(.a(dm_int_st5_29[3]), .b(dm_int_st5_29[4]), .cin(dm_int_st5_29[5]), .s(dm_int_st6_29[3]), .cout(dm_int_st6_30[1]));
	// Bit 30
	full_adder FA724(.a(dm_int_st5_30[0]), .b(dm_int_st5_30[1]), .cin(dm_int_st5_30[2]), .s(dm_int_st6_30[2]), .cout(dm_int_st6_31[0]));
	full_adder FA725(.a(dm_int_st5_30[3]), .b(dm_int_st5_30[4]), .cin(dm_int_st5_30[5]), .s(dm_int_st6_30[3]), .cout(dm_int_st6_31[1]));
	// Bit 31
	full_adder FA726(.a(dm_int_st5_31[0]), .b(dm_int_st5_31[1]), .cin(dm_int_st5_31[2]), .s(dm_int_st6_31[2]), .cout(dm_int_st6_32[0]));
	full_adder FA727(.a(dm_int_st5_31[3]), .b(dm_int_st5_31[4]), .cin(dm_int_st5_31[5]), .s(dm_int_st6_31[3]), .cout(dm_int_st6_32[1]));
	// Bit 32
	full_adder FA728(.a(dm_int_st5_32[0]), .b(dm_int_st5_32[1]), .cin(dm_int_st5_32[2]), .s(dm_int_st6_32[2]), .cout(dm_int_st6_33[0]));
	full_adder FA729(.a(dm_int_st5_32[3]), .b(dm_int_st5_32[4]), .cin(dm_int_st5_32[5]), .s(dm_int_st6_32[3]), .cout(dm_int_st6_33[1]));
	// Bit 33
	full_adder FA730(.a(dm_int_st5_33[0]), .b(dm_int_st5_33[1]), .cin(dm_int_st5_33[2]), .s(dm_int_st6_33[2]), .cout(dm_int_st6_34[0]));
	full_adder FA731(.a(dm_int_st5_33[3]), .b(dm_int_st5_33[4]), .cin(dm_int_st5_33[5]), .s(dm_int_st6_33[3]), .cout(dm_int_st6_34[1]));
	// Bit 34
	full_adder FA732(.a(dm_int_st5_34[0]), .b(dm_int_st5_34[1]), .cin(dm_int_st5_34[2]), .s(dm_int_st6_34[2]), .cout(dm_int_st6_35[0]));
	full_adder FA733(.a(dm_int_st5_34[3]), .b(dm_int_st5_34[4]), .cin(dm_int_st5_34[5]), .s(dm_int_st6_34[3]), .cout(dm_int_st6_35[1]));
	// Bit 35
	full_adder FA734(.a(dm_int_st5_35[0]), .b(dm_int_st5_35[1]), .cin(dm_int_st5_35[2]), .s(dm_int_st6_35[2]), .cout(dm_int_st6_36[0]));
	full_adder FA735(.a(dm_int_st5_35[3]), .b(dm_int_st5_35[4]), .cin(dm_int_st5_35[5]), .s(dm_int_st6_35[3]), .cout(dm_int_st6_36[1]));
	// Bit 36
	full_adder FA736(.a(dm_int_st5_36[0]), .b(dm_int_st5_36[1]), .cin(dm_int_st5_36[2]), .s(dm_int_st6_36[2]), .cout(dm_int_st6_37[0]));
	full_adder FA737(.a(dm_int_st5_36[3]), .b(dm_int_st5_36[4]), .cin(dm_int_st5_36[5]), .s(dm_int_st6_36[3]), .cout(dm_int_st6_37[1]));
	// Bit 37
	full_adder FA738(.a(dm_int_st5_37[0]), .b(dm_int_st5_37[1]), .cin(dm_int_st5_37[2]), .s(dm_int_st6_37[2]), .cout(dm_int_st6_38[0]));
	full_adder FA739(.a(dm_int_st5_37[3]), .b(dm_int_st5_37[4]), .cin(dm_int_st5_37[5]), .s(dm_int_st6_37[3]), .cout(dm_int_st6_38[1]));
	// Bit 38
	full_adder FA740(.a(dm_int_st5_38[0]), .b(dm_int_st5_38[1]), .cin(dm_int_st5_38[2]), .s(dm_int_st6_38[2]), .cout(dm_int_st6_39[0]));
	full_adder FA741(.a(dm_int_st5_38[3]), .b(dm_int_st5_38[4]), .cin(dm_int_st5_38[5]), .s(dm_int_st6_38[3]), .cout(dm_int_st6_39[1]));
	// Bit 39
	full_adder FA742(.a(dm_int_st5_39[0]), .b(dm_int_st5_39[1]), .cin(dm_int_st5_39[2]), .s(dm_int_st6_39[2]), .cout(dm_int_st6_40[0]));
	full_adder FA743(.a(dm_int_st5_39[3]), .b(dm_int_st5_39[4]), .cin(dm_int_st5_39[5]), .s(dm_int_st6_39[3]), .cout(dm_int_st6_40[1]));
	// Bit 40
	full_adder FA744(.a(dm_int_st5_40[0]), .b(dm_int_st5_40[1]), .cin(dm_int_st5_40[2]), .s(dm_int_st6_40[2]), .cout(dm_int_st6_41[0]));
	full_adder FA745(.a(dm_int_st5_40[3]), .b(dm_int_st5_40[4]), .cin(dm_int_st5_40[5]), .s(dm_int_st6_40[3]), .cout(dm_int_st6_41[1]));
	// Bit 41
	full_adder FA746(.a(dm_int_st5_41[0]), .b(dm_int_st5_41[1]), .cin(dm_int_st5_41[2]), .s(dm_int_st6_41[2]), .cout(dm_int_st6_42[0]));
	full_adder FA747(.a(dm_int_st5_41[3]), .b(dm_int_st5_41[4]), .cin(dm_int_st5_41[5]), .s(dm_int_st6_41[3]), .cout(dm_int_st6_42[1]));
	// Bit 42
	full_adder FA748(.a(dm_int_st5_42[0]), .b(dm_int_st5_42[1]), .cin(dm_int_st5_42[2]), .s(dm_int_st6_42[2]), .cout(dm_int_st6_43[0]));
	full_adder FA749(.a(dm_int_st5_42[3]), .b(dm_int_st5_42[4]), .cin(dm_int_st5_42[5]), .s(dm_int_st6_42[3]), .cout(dm_int_st6_43[1]));
	// Bit 43
	full_adder FA750(.a(dm_int_st5_43[0]), .b(dm_int_st5_43[1]), .cin(dm_int_st5_43[2]), .s(dm_int_st6_43[2]), .cout(dm_int_st6_44[0]));
	full_adder FA751(.a(dm_int_st5_43[3]), .b(dm_int_st5_43[4]), .cin(dm_int_st5_43[5]), .s(dm_int_st6_43[3]), .cout(dm_int_st6_44[1]));
	// Bit 44
	full_adder FA752(.a(dm_int_st5_44[0]), .b(dm_int_st5_44[1]), .cin(dm_int_st5_44[2]), .s(dm_int_st6_44[2]), .cout(dm_int_st6_45[0]));
	full_adder FA753(.a(dm_int_st5_44[3]), .b(dm_int_st5_44[4]), .cin(dm_int_st5_44[5]), .s(dm_int_st6_44[3]), .cout(dm_int_st6_45[1]));
	// Bit 45
	full_adder FA754(.a(dm_int_st5_45[0]), .b(dm_int_st5_45[1]), .cin(dm_int_st5_45[2]), .s(dm_int_st6_45[2]), .cout(dm_int_st6_46[0]));
	full_adder FA755(.a(dm_int_st5_45[3]), .b(dm_int_st5_45[4]), .cin(dm_int_st5_45[5]), .s(dm_int_st6_45[3]), .cout(dm_int_st6_46[1]));
	// Bit 46
	full_adder FA756(.a(dm_int_st5_46[0]), .b(dm_int_st5_46[1]), .cin(dm_int_st5_46[2]), .s(dm_int_st6_46[2]), .cout(dm_int_st6_47[0]));
	full_adder FA757(.a(dm_int_st5_46[3]), .b(dm_int_st5_46[4]), .cin(dm_int_st5_46[5]), .s(dm_int_st6_46[3]), .cout(dm_int_st6_47[1]));
	// Bit 47
	full_adder FA758(.a(dm_int_st5_47[0]), .b(dm_int_st5_47[1]), .cin(dm_int_st5_47[2]), .s(dm_int_st6_47[2]), .cout(dm_int_st6_48[0]));
	full_adder FA759(.a(dm_int_st5_47[3]), .b(dm_int_st5_47[4]), .cin(dm_int_st5_47[5]), .s(dm_int_st6_47[3]), .cout(dm_int_st6_48[1]));
	// Bit 48
	full_adder FA760(.a(dm_int_st5_48[0]), .b(dm_int_st5_48[1]), .cin(dm_int_st5_48[2]), .s(dm_int_st6_48[2]), .cout(dm_int_st6_49[0]));
	full_adder FA761(.a(dm_int_st5_48[3]), .b(dm_int_st5_48[4]), .cin(dm_int_st5_48[5]), .s(dm_int_st6_48[3]), .cout(dm_int_st6_49[1]));
	// Bit 49
	full_adder FA762(.a(dm_int_st5_49[0]), .b(dm_int_st5_49[1]), .cin(dm_int_st5_49[2]), .s(dm_int_st6_49[2]), .cout(dm_int_st6_50[0]));
	full_adder FA763(.a(dm_int_st5_49[3]), .b(dm_int_st5_49[4]), .cin(dm_int_st5_49[5]), .s(dm_int_st6_49[3]), .cout(dm_int_st6_50[1]));
	// Bit 50
	full_adder FA764(.a(dm_int_st5_50[0]), .b(dm_int_st5_50[1]), .cin(dm_int_st5_50[2]), .s(dm_int_st6_50[2]), .cout(dm_int_st6_51[0]));
	full_adder FA765(.a(dm_int_st5_50[3]), .b(dm_int_st5_50[4]), .cin(dm_int_st5_50[5]), .s(dm_int_st6_50[3]), .cout(dm_int_st6_51[1]));
	// Bit 51
	full_adder FA766(.a(dm_int_st5_51[0]), .b(dm_int_st5_51[1]), .cin(dm_int_st5_51[2]), .s(dm_int_st6_51[2]), .cout(dm_int_st6_52[0]));
	full_adder FA767(.a(dm_int_st5_51[3]), .b(dm_int_st5_51[4]), .cin(dm_int_st5_51[5]), .s(dm_int_st6_51[3]), .cout(dm_int_st6_52[1]));
	// Bit 52
	full_adder FA768(.a(dm_int_st5_52[0]), .b(dm_int_st5_52[1]), .cin(dm_int_st5_52[2]), .s(dm_int_st6_52[2]), .cout(dm_int_st6_53[0]));
	full_adder FA769(.a(dm_int_st5_52[3]), .b(dm_int_st5_52[4]), .cin(dm_int_st5_52[5]), .s(dm_int_st6_52[3]), .cout(dm_int_st6_53[1]));
	// Bit 53
	full_adder FA770(.a(dm_int_st5_53[0]), .b(dm_int_st5_53[1]), .cin(dm_int_st5_53[2]), .s(dm_int_st6_53[2]), .cout(dm_int_st6_54[0]));
	full_adder FA771(.a(dm_int_st5_53[3]), .b(dm_int_st5_53[4]), .cin(dm_int_st5_53[5]), .s(dm_int_st6_53[3]), .cout(dm_int_st6_54[1]));
	// Bit 54
	full_adder FA772(.a(dm_int_st5_54[0]), .b(dm_int_st5_54[1]), .cin(dm_int_st5_54[2]), .s(dm_int_st6_54[2]), .cout(dm_int_st6_55[0]));
	full_adder FA773(.a(dm_int_st5_54[3]), .b(dm_int_st5_54[4]), .cin(dm_int_st5_54[5]), .s(dm_int_st6_54[3]), .cout(dm_int_st6_55[1]));
	// Bit 55
	full_adder FA774(.a(dm_int_st5_55[0]), .b(dm_int_st5_55[1]), .cin(dm_int_st5_55[2]), .s(dm_int_st6_55[2]), .cout(dm_int_st6_56[0]));
	full_adder FA775(.a(dm_int_st5_55[3]), .b(dm_int_st5_55[4]), .cin(dm_int_st5_55[5]), .s(dm_int_st6_55[3]), .cout(dm_int_st6_56[1]));
	// Bit 56
	full_adder FA776(.a(dm_int_st5_56[0]), .b(dm_int_st5_56[1]), .cin(dm_int_st5_56[2]), .s(dm_int_st6_56[2]), .cout(dm_int_st6_57[0]));
	full_adder FA777(.a(dm_int_st5_56[3]), .b(dm_int_st5_56[4]), .cin(dm_int_st5_56[5]), .s(dm_int_st6_56[3]), .cout(dm_int_st6_57[1]));
	// Bit 57
	full_adder FA778(.a(dm_int_st5_57[0]), .b(dm_int_st5_57[1]), .cin(dm_int_st5_57[2]), .s(dm_int_st6_57[2]), .cout(dm_int_st6_58[0]));
	full_adder FA779(.a(dm_int_st5_57[3]), .b(dm_int_st5_57[4]), .cin(dm_int_st5_57[5]), .s(dm_int_st6_57[3]), .cout(dm_int_st6_58[1]));
	// Bit 58
	full_adder FA780(.a(dm_int_st5_58[0]), .b(dm_int_st5_58[1]), .cin(dm_int_st5_58[2]), .s(dm_int_st6_58[2]), .cout(dm_int_st6_59[0]));
	full_adder FA781(.a(dm_int_st5_58[3]), .b(dm_int_st5_58[4]), .cin(dm_int_st5_58[5]), .s(dm_int_st6_58[3]), .cout(dm_int_st6_59[1]));
	// Bit 59
	full_adder FA782(.a(dm_int_st5_59[0]), .b(dm_int_st5_59[1]), .cin(dm_int_st5_59[2]), .s(dm_int_st6_59[2]), .cout(dm_int_st6_60[0]));
	assign dm_int_st6_59[3] = dm_int_st5_59[3];
	// Bit 60
	assign dm_int_st6_60[1] = dm_int_st5_60[0];
	assign dm_int_st6_60[2] = dm_int_st5_60[1];
	assign dm_int_st6_60[3] = dm_int_st5_60[2];
	// Bit 61
	assign dm_int_st6_61[0] = dm_int_st5_61[0];
	assign dm_int_st6_61[1] = dm_int_st5_61[1];
	// Bit 62
	assign dm_int_st6_62[0] = dm_int_st5_62[0];

	//// Stage 7 ////
	wire [0:0] dm_int_st7_0;
	wire [1:0] dm_int_st7_1;
	wire [2:0] dm_int_st7_2;
	wire [2:0] dm_int_st7_3;
	wire [2:0] dm_int_st7_4;
	wire [2:0] dm_int_st7_5;
	wire [2:0] dm_int_st7_6;
	wire [2:0] dm_int_st7_7;
	wire [2:0] dm_int_st7_8;
	wire [2:0] dm_int_st7_9;
	wire [2:0] dm_int_st7_10;
	wire [2:0] dm_int_st7_11;
	wire [2:0] dm_int_st7_12;
	wire [2:0] dm_int_st7_13;
	wire [2:0] dm_int_st7_14;
	wire [2:0] dm_int_st7_15;
	wire [2:0] dm_int_st7_16;
	wire [2:0] dm_int_st7_17;
	wire [2:0] dm_int_st7_18;
	wire [2:0] dm_int_st7_19;
	wire [2:0] dm_int_st7_20;
	wire [2:0] dm_int_st7_21;
	wire [2:0] dm_int_st7_22;
	wire [2:0] dm_int_st7_23;
	wire [2:0] dm_int_st7_24;
	wire [2:0] dm_int_st7_25;
	wire [2:0] dm_int_st7_26;
	wire [2:0] dm_int_st7_27;
	wire [2:0] dm_int_st7_28;
	wire [2:0] dm_int_st7_29;
	wire [2:0] dm_int_st7_30;
	wire [2:0] dm_int_st7_31;
	wire [2:0] dm_int_st7_32;
	wire [2:0] dm_int_st7_33;
	wire [2:0] dm_int_st7_34;
	wire [2:0] dm_int_st7_35;
	wire [2:0] dm_int_st7_36;
	wire [2:0] dm_int_st7_37;
	wire [2:0] dm_int_st7_38;
	wire [2:0] dm_int_st7_39;
	wire [2:0] dm_int_st7_40;
	wire [2:0] dm_int_st7_41;
	wire [2:0] dm_int_st7_42;
	wire [2:0] dm_int_st7_43;
	wire [2:0] dm_int_st7_44;
	wire [2:0] dm_int_st7_45;
	wire [2:0] dm_int_st7_46;
	wire [2:0] dm_int_st7_47;
	wire [2:0] dm_int_st7_48;
	wire [2:0] dm_int_st7_49;
	wire [2:0] dm_int_st7_50;
	wire [2:0] dm_int_st7_51;
	wire [2:0] dm_int_st7_52;
	wire [2:0] dm_int_st7_53;
	wire [2:0] dm_int_st7_54;
	wire [2:0] dm_int_st7_55;
	wire [2:0] dm_int_st7_56;
	wire [2:0] dm_int_st7_57;
	wire [2:0] dm_int_st7_58;
	wire [2:0] dm_int_st7_59;
	wire [2:0] dm_int_st7_60;
	wire [2:0] dm_int_st7_61;
	wire [0:0] dm_int_st7_62;

	// Bit 0
	assign dm_int_st7_0[0] = dm_int_st6_0[0];
	// Bit 1
	assign dm_int_st7_1[0] = dm_int_st6_1[0];
	assign dm_int_st7_1[1] = dm_int_st6_1[1];
	// Bit 2
	assign dm_int_st7_2[0] = dm_int_st6_2[0];
	assign dm_int_st7_2[1] = dm_int_st6_2[1];
	assign dm_int_st7_2[2] = dm_int_st6_2[2];
	// Bit 3
	half_adder HA29(.a(dm_int_st6_3[0]), .b(dm_int_st6_3[1]), .s(dm_int_st7_3[0]), .cout(dm_int_st7_4[0]));
	assign dm_int_st7_3[1] = dm_int_st6_3[2];
	assign dm_int_st7_3[2] = dm_int_st6_3[3];
	// Bit 4
	full_adder FA783(.a(dm_int_st6_4[0]), .b(dm_int_st6_4[1]), .cin(dm_int_st6_4[2]), .s(dm_int_st7_4[1]), .cout(dm_int_st7_5[0]));
	assign dm_int_st7_4[2] = dm_int_st6_4[3];
	// Bit 5
	full_adder FA784(.a(dm_int_st6_5[0]), .b(dm_int_st6_5[1]), .cin(dm_int_st6_5[2]), .s(dm_int_st7_5[1]), .cout(dm_int_st7_6[0]));
	assign dm_int_st7_5[2] = dm_int_st6_5[3];
	// Bit 6
	full_adder FA785(.a(dm_int_st6_6[0]), .b(dm_int_st6_6[1]), .cin(dm_int_st6_6[2]), .s(dm_int_st7_6[1]), .cout(dm_int_st7_7[0]));
	assign dm_int_st7_6[2] = dm_int_st6_6[3];
	// Bit 7
	full_adder FA786(.a(dm_int_st6_7[0]), .b(dm_int_st6_7[1]), .cin(dm_int_st6_7[2]), .s(dm_int_st7_7[1]), .cout(dm_int_st7_8[0]));
	assign dm_int_st7_7[2] = dm_int_st6_7[3];
	// Bit 8
	full_adder FA787(.a(dm_int_st6_8[0]), .b(dm_int_st6_8[1]), .cin(dm_int_st6_8[2]), .s(dm_int_st7_8[1]), .cout(dm_int_st7_9[0]));
	assign dm_int_st7_8[2] = dm_int_st6_8[3];
	// Bit 9
	full_adder FA788(.a(dm_int_st6_9[0]), .b(dm_int_st6_9[1]), .cin(dm_int_st6_9[2]), .s(dm_int_st7_9[1]), .cout(dm_int_st7_10[0]));
	assign dm_int_st7_9[2] = dm_int_st6_9[3];
	// Bit 10
	full_adder FA789(.a(dm_int_st6_10[0]), .b(dm_int_st6_10[1]), .cin(dm_int_st6_10[2]), .s(dm_int_st7_10[1]), .cout(dm_int_st7_11[0]));
	assign dm_int_st7_10[2] = dm_int_st6_10[3];
	// Bit 11
	full_adder FA790(.a(dm_int_st6_11[0]), .b(dm_int_st6_11[1]), .cin(dm_int_st6_11[2]), .s(dm_int_st7_11[1]), .cout(dm_int_st7_12[0]));
	assign dm_int_st7_11[2] = dm_int_st6_11[3];
	// Bit 12
	full_adder FA791(.a(dm_int_st6_12[0]), .b(dm_int_st6_12[1]), .cin(dm_int_st6_12[2]), .s(dm_int_st7_12[1]), .cout(dm_int_st7_13[0]));
	assign dm_int_st7_12[2] = dm_int_st6_12[3];
	// Bit 13
	full_adder FA792(.a(dm_int_st6_13[0]), .b(dm_int_st6_13[1]), .cin(dm_int_st6_13[2]), .s(dm_int_st7_13[1]), .cout(dm_int_st7_14[0]));
	assign dm_int_st7_13[2] = dm_int_st6_13[3];
	// Bit 14
	full_adder FA793(.a(dm_int_st6_14[0]), .b(dm_int_st6_14[1]), .cin(dm_int_st6_14[2]), .s(dm_int_st7_14[1]), .cout(dm_int_st7_15[0]));
	assign dm_int_st7_14[2] = dm_int_st6_14[3];
	// Bit 15
	full_adder FA794(.a(dm_int_st6_15[0]), .b(dm_int_st6_15[1]), .cin(dm_int_st6_15[2]), .s(dm_int_st7_15[1]), .cout(dm_int_st7_16[0]));
	assign dm_int_st7_15[2] = dm_int_st6_15[3];
	// Bit 16
	full_adder FA795(.a(dm_int_st6_16[0]), .b(dm_int_st6_16[1]), .cin(dm_int_st6_16[2]), .s(dm_int_st7_16[1]), .cout(dm_int_st7_17[0]));
	assign dm_int_st7_16[2] = dm_int_st6_16[3];
	// Bit 17
	full_adder FA796(.a(dm_int_st6_17[0]), .b(dm_int_st6_17[1]), .cin(dm_int_st6_17[2]), .s(dm_int_st7_17[1]), .cout(dm_int_st7_18[0]));
	assign dm_int_st7_17[2] = dm_int_st6_17[3];
	// Bit 18
	full_adder FA797(.a(dm_int_st6_18[0]), .b(dm_int_st6_18[1]), .cin(dm_int_st6_18[2]), .s(dm_int_st7_18[1]), .cout(dm_int_st7_19[0]));
	assign dm_int_st7_18[2] = dm_int_st6_18[3];
	// Bit 19
	full_adder FA798(.a(dm_int_st6_19[0]), .b(dm_int_st6_19[1]), .cin(dm_int_st6_19[2]), .s(dm_int_st7_19[1]), .cout(dm_int_st7_20[0]));
	assign dm_int_st7_19[2] = dm_int_st6_19[3];
	// Bit 20
	full_adder FA799(.a(dm_int_st6_20[0]), .b(dm_int_st6_20[1]), .cin(dm_int_st6_20[2]), .s(dm_int_st7_20[1]), .cout(dm_int_st7_21[0]));
	assign dm_int_st7_20[2] = dm_int_st6_20[3];
	// Bit 21
	full_adder FA800(.a(dm_int_st6_21[0]), .b(dm_int_st6_21[1]), .cin(dm_int_st6_21[2]), .s(dm_int_st7_21[1]), .cout(dm_int_st7_22[0]));
	assign dm_int_st7_21[2] = dm_int_st6_21[3];
	// Bit 22
	full_adder FA801(.a(dm_int_st6_22[0]), .b(dm_int_st6_22[1]), .cin(dm_int_st6_22[2]), .s(dm_int_st7_22[1]), .cout(dm_int_st7_23[0]));
	assign dm_int_st7_22[2] = dm_int_st6_22[3];
	// Bit 23
	full_adder FA802(.a(dm_int_st6_23[0]), .b(dm_int_st6_23[1]), .cin(dm_int_st6_23[2]), .s(dm_int_st7_23[1]), .cout(dm_int_st7_24[0]));
	assign dm_int_st7_23[2] = dm_int_st6_23[3];
	// Bit 24
	full_adder FA803(.a(dm_int_st6_24[0]), .b(dm_int_st6_24[1]), .cin(dm_int_st6_24[2]), .s(dm_int_st7_24[1]), .cout(dm_int_st7_25[0]));
	assign dm_int_st7_24[2] = dm_int_st6_24[3];
	// Bit 25
	full_adder FA804(.a(dm_int_st6_25[0]), .b(dm_int_st6_25[1]), .cin(dm_int_st6_25[2]), .s(dm_int_st7_25[1]), .cout(dm_int_st7_26[0]));
	assign dm_int_st7_25[2] = dm_int_st6_25[3];
	// Bit 26
	full_adder FA805(.a(dm_int_st6_26[0]), .b(dm_int_st6_26[1]), .cin(dm_int_st6_26[2]), .s(dm_int_st7_26[1]), .cout(dm_int_st7_27[0]));
	assign dm_int_st7_26[2] = dm_int_st6_26[3];
	// Bit 27
	full_adder FA806(.a(dm_int_st6_27[0]), .b(dm_int_st6_27[1]), .cin(dm_int_st6_27[2]), .s(dm_int_st7_27[1]), .cout(dm_int_st7_28[0]));
	assign dm_int_st7_27[2] = dm_int_st6_27[3];
	// Bit 28
	full_adder FA807(.a(dm_int_st6_28[0]), .b(dm_int_st6_28[1]), .cin(dm_int_st6_28[2]), .s(dm_int_st7_28[1]), .cout(dm_int_st7_29[0]));
	assign dm_int_st7_28[2] = dm_int_st6_28[3];
	// Bit 29
	full_adder FA808(.a(dm_int_st6_29[0]), .b(dm_int_st6_29[1]), .cin(dm_int_st6_29[2]), .s(dm_int_st7_29[1]), .cout(dm_int_st7_30[0]));
	assign dm_int_st7_29[2] = dm_int_st6_29[3];
	// Bit 30
	full_adder FA809(.a(dm_int_st6_30[0]), .b(dm_int_st6_30[1]), .cin(dm_int_st6_30[2]), .s(dm_int_st7_30[1]), .cout(dm_int_st7_31[0]));
	assign dm_int_st7_30[2] = dm_int_st6_30[3];
	// Bit 31
	full_adder FA810(.a(dm_int_st6_31[0]), .b(dm_int_st6_31[1]), .cin(dm_int_st6_31[2]), .s(dm_int_st7_31[1]), .cout(dm_int_st7_32[0]));
	assign dm_int_st7_31[2] = dm_int_st6_31[3];
	// Bit 32
	full_adder FA811(.a(dm_int_st6_32[0]), .b(dm_int_st6_32[1]), .cin(dm_int_st6_32[2]), .s(dm_int_st7_32[1]), .cout(dm_int_st7_33[0]));
	assign dm_int_st7_32[2] = dm_int_st6_32[3];
	// Bit 33
	full_adder FA812(.a(dm_int_st6_33[0]), .b(dm_int_st6_33[1]), .cin(dm_int_st6_33[2]), .s(dm_int_st7_33[1]), .cout(dm_int_st7_34[0]));
	assign dm_int_st7_33[2] = dm_int_st6_33[3];
	// Bit 34
	full_adder FA813(.a(dm_int_st6_34[0]), .b(dm_int_st6_34[1]), .cin(dm_int_st6_34[2]), .s(dm_int_st7_34[1]), .cout(dm_int_st7_35[0]));
	assign dm_int_st7_34[2] = dm_int_st6_34[3];
	// Bit 35
	full_adder FA814(.a(dm_int_st6_35[0]), .b(dm_int_st6_35[1]), .cin(dm_int_st6_35[2]), .s(dm_int_st7_35[1]), .cout(dm_int_st7_36[0]));
	assign dm_int_st7_35[2] = dm_int_st6_35[3];
	// Bit 36
	full_adder FA815(.a(dm_int_st6_36[0]), .b(dm_int_st6_36[1]), .cin(dm_int_st6_36[2]), .s(dm_int_st7_36[1]), .cout(dm_int_st7_37[0]));
	assign dm_int_st7_36[2] = dm_int_st6_36[3];
	// Bit 37
	full_adder FA816(.a(dm_int_st6_37[0]), .b(dm_int_st6_37[1]), .cin(dm_int_st6_37[2]), .s(dm_int_st7_37[1]), .cout(dm_int_st7_38[0]));
	assign dm_int_st7_37[2] = dm_int_st6_37[3];
	// Bit 38
	full_adder FA817(.a(dm_int_st6_38[0]), .b(dm_int_st6_38[1]), .cin(dm_int_st6_38[2]), .s(dm_int_st7_38[1]), .cout(dm_int_st7_39[0]));
	assign dm_int_st7_38[2] = dm_int_st6_38[3];
	// Bit 39
	full_adder FA818(.a(dm_int_st6_39[0]), .b(dm_int_st6_39[1]), .cin(dm_int_st6_39[2]), .s(dm_int_st7_39[1]), .cout(dm_int_st7_40[0]));
	assign dm_int_st7_39[2] = dm_int_st6_39[3];
	// Bit 40
	full_adder FA819(.a(dm_int_st6_40[0]), .b(dm_int_st6_40[1]), .cin(dm_int_st6_40[2]), .s(dm_int_st7_40[1]), .cout(dm_int_st7_41[0]));
	assign dm_int_st7_40[2] = dm_int_st6_40[3];
	// Bit 41
	full_adder FA820(.a(dm_int_st6_41[0]), .b(dm_int_st6_41[1]), .cin(dm_int_st6_41[2]), .s(dm_int_st7_41[1]), .cout(dm_int_st7_42[0]));
	assign dm_int_st7_41[2] = dm_int_st6_41[3];
	// Bit 42
	full_adder FA821(.a(dm_int_st6_42[0]), .b(dm_int_st6_42[1]), .cin(dm_int_st6_42[2]), .s(dm_int_st7_42[1]), .cout(dm_int_st7_43[0]));
	assign dm_int_st7_42[2] = dm_int_st6_42[3];
	// Bit 43
	full_adder FA822(.a(dm_int_st6_43[0]), .b(dm_int_st6_43[1]), .cin(dm_int_st6_43[2]), .s(dm_int_st7_43[1]), .cout(dm_int_st7_44[0]));
	assign dm_int_st7_43[2] = dm_int_st6_43[3];
	// Bit 44
	full_adder FA823(.a(dm_int_st6_44[0]), .b(dm_int_st6_44[1]), .cin(dm_int_st6_44[2]), .s(dm_int_st7_44[1]), .cout(dm_int_st7_45[0]));
	assign dm_int_st7_44[2] = dm_int_st6_44[3];
	// Bit 45
	full_adder FA824(.a(dm_int_st6_45[0]), .b(dm_int_st6_45[1]), .cin(dm_int_st6_45[2]), .s(dm_int_st7_45[1]), .cout(dm_int_st7_46[0]));
	assign dm_int_st7_45[2] = dm_int_st6_45[3];
	// Bit 46
	full_adder FA825(.a(dm_int_st6_46[0]), .b(dm_int_st6_46[1]), .cin(dm_int_st6_46[2]), .s(dm_int_st7_46[1]), .cout(dm_int_st7_47[0]));
	assign dm_int_st7_46[2] = dm_int_st6_46[3];
	// Bit 47
	full_adder FA826(.a(dm_int_st6_47[0]), .b(dm_int_st6_47[1]), .cin(dm_int_st6_47[2]), .s(dm_int_st7_47[1]), .cout(dm_int_st7_48[0]));
	assign dm_int_st7_47[2] = dm_int_st6_47[3];
	// Bit 48
	full_adder FA827(.a(dm_int_st6_48[0]), .b(dm_int_st6_48[1]), .cin(dm_int_st6_48[2]), .s(dm_int_st7_48[1]), .cout(dm_int_st7_49[0]));
	assign dm_int_st7_48[2] = dm_int_st6_48[3];
	// Bit 49
	full_adder FA828(.a(dm_int_st6_49[0]), .b(dm_int_st6_49[1]), .cin(dm_int_st6_49[2]), .s(dm_int_st7_49[1]), .cout(dm_int_st7_50[0]));
	assign dm_int_st7_49[2] = dm_int_st6_49[3];
	// Bit 50
	full_adder FA829(.a(dm_int_st6_50[0]), .b(dm_int_st6_50[1]), .cin(dm_int_st6_50[2]), .s(dm_int_st7_50[1]), .cout(dm_int_st7_51[0]));
	assign dm_int_st7_50[2] = dm_int_st6_50[3];
	// Bit 51
	full_adder FA830(.a(dm_int_st6_51[0]), .b(dm_int_st6_51[1]), .cin(dm_int_st6_51[2]), .s(dm_int_st7_51[1]), .cout(dm_int_st7_52[0]));
	assign dm_int_st7_51[2] = dm_int_st6_51[3];
	// Bit 52
	full_adder FA831(.a(dm_int_st6_52[0]), .b(dm_int_st6_52[1]), .cin(dm_int_st6_52[2]), .s(dm_int_st7_52[1]), .cout(dm_int_st7_53[0]));
	assign dm_int_st7_52[2] = dm_int_st6_52[3];
	// Bit 53
	full_adder FA832(.a(dm_int_st6_53[0]), .b(dm_int_st6_53[1]), .cin(dm_int_st6_53[2]), .s(dm_int_st7_53[1]), .cout(dm_int_st7_54[0]));
	assign dm_int_st7_53[2] = dm_int_st6_53[3];
	// Bit 54
	full_adder FA833(.a(dm_int_st6_54[0]), .b(dm_int_st6_54[1]), .cin(dm_int_st6_54[2]), .s(dm_int_st7_54[1]), .cout(dm_int_st7_55[0]));
	assign dm_int_st7_54[2] = dm_int_st6_54[3];
	// Bit 55
	full_adder FA834(.a(dm_int_st6_55[0]), .b(dm_int_st6_55[1]), .cin(dm_int_st6_55[2]), .s(dm_int_st7_55[1]), .cout(dm_int_st7_56[0]));
	assign dm_int_st7_55[2] = dm_int_st6_55[3];
	// Bit 56
	full_adder FA835(.a(dm_int_st6_56[0]), .b(dm_int_st6_56[1]), .cin(dm_int_st6_56[2]), .s(dm_int_st7_56[1]), .cout(dm_int_st7_57[0]));
	assign dm_int_st7_56[2] = dm_int_st6_56[3];
	// Bit 57
	full_adder FA836(.a(dm_int_st6_57[0]), .b(dm_int_st6_57[1]), .cin(dm_int_st6_57[2]), .s(dm_int_st7_57[1]), .cout(dm_int_st7_58[0]));
	assign dm_int_st7_57[2] = dm_int_st6_57[3];
	// Bit 58
	full_adder FA837(.a(dm_int_st6_58[0]), .b(dm_int_st6_58[1]), .cin(dm_int_st6_58[2]), .s(dm_int_st7_58[1]), .cout(dm_int_st7_59[0]));
	assign dm_int_st7_58[2] = dm_int_st6_58[3];
	// Bit 59
	full_adder FA838(.a(dm_int_st6_59[0]), .b(dm_int_st6_59[1]), .cin(dm_int_st6_59[2]), .s(dm_int_st7_59[1]), .cout(dm_int_st7_60[0]));
	assign dm_int_st7_59[2] = dm_int_st6_59[3];
	// Bit 60
	full_adder FA839(.a(dm_int_st6_60[0]), .b(dm_int_st6_60[1]), .cin(dm_int_st6_60[2]), .s(dm_int_st7_60[1]), .cout(dm_int_st7_61[0]));
	assign dm_int_st7_60[2] = dm_int_st6_60[3];
	// Bit 61
	assign dm_int_st7_61[1] = dm_int_st6_61[0];
	assign dm_int_st7_61[2] = dm_int_st6_61[1];
	// Bit 62
	assign dm_int_st7_62[0] = dm_int_st6_62[0];

	//// Stage 8 ////
	wire [0:0] dm_int_st8_0;
	wire [1:0] dm_int_st8_1;
	wire [1:0] dm_int_st8_2;
	wire [1:0] dm_int_st8_3;
	wire [1:0] dm_int_st8_4;
	wire [1:0] dm_int_st8_5;
	wire [1:0] dm_int_st8_6;
	wire [1:0] dm_int_st8_7;
	wire [1:0] dm_int_st8_8;
	wire [1:0] dm_int_st8_9;
	wire [1:0] dm_int_st8_10;
	wire [1:0] dm_int_st8_11;
	wire [1:0] dm_int_st8_12;
	wire [1:0] dm_int_st8_13;
	wire [1:0] dm_int_st8_14;
	wire [1:0] dm_int_st8_15;
	wire [1:0] dm_int_st8_16;
	wire [1:0] dm_int_st8_17;
	wire [1:0] dm_int_st8_18;
	wire [1:0] dm_int_st8_19;
	wire [1:0] dm_int_st8_20;
	wire [1:0] dm_int_st8_21;
	wire [1:0] dm_int_st8_22;
	wire [1:0] dm_int_st8_23;
	wire [1:0] dm_int_st8_24;
	wire [1:0] dm_int_st8_25;
	wire [1:0] dm_int_st8_26;
	wire [1:0] dm_int_st8_27;
	wire [1:0] dm_int_st8_28;
	wire [1:0] dm_int_st8_29;
	wire [1:0] dm_int_st8_30;
	wire [1:0] dm_int_st8_31;
	wire [1:0] dm_int_st8_32;
	wire [1:0] dm_int_st8_33;
	wire [1:0] dm_int_st8_34;
	wire [1:0] dm_int_st8_35;
	wire [1:0] dm_int_st8_36;
	wire [1:0] dm_int_st8_37;
	wire [1:0] dm_int_st8_38;
	wire [1:0] dm_int_st8_39;
	wire [1:0] dm_int_st8_40;
	wire [1:0] dm_int_st8_41;
	wire [1:0] dm_int_st8_42;
	wire [1:0] dm_int_st8_43;
	wire [1:0] dm_int_st8_44;
	wire [1:0] dm_int_st8_45;
	wire [1:0] dm_int_st8_46;
	wire [1:0] dm_int_st8_47;
	wire [1:0] dm_int_st8_48;
	wire [1:0] dm_int_st8_49;
	wire [1:0] dm_int_st8_50;
	wire [1:0] dm_int_st8_51;
	wire [1:0] dm_int_st8_52;
	wire [1:0] dm_int_st8_53;
	wire [1:0] dm_int_st8_54;
	wire [1:0] dm_int_st8_55;
	wire [1:0] dm_int_st8_56;
	wire [1:0] dm_int_st8_57;
	wire [1:0] dm_int_st8_58;
	wire [1:0] dm_int_st8_59;
	wire [1:0] dm_int_st8_60;
	wire [1:0] dm_int_st8_61;
	wire [1:0] dm_int_st8_62;

	// Bit 0
	assign dm_int_st8_0[0] = dm_int_st7_0[0];
	// Bit 1
	assign dm_int_st8_1[0] = dm_int_st7_1[0];
	assign dm_int_st8_1[1] = dm_int_st7_1[1];
	// Bit 2
	half_adder HA30(.a(dm_int_st7_2[0]), .b(dm_int_st7_2[1]), .s(dm_int_st8_2[0]), .cout(dm_int_st8_3[0]));
	assign dm_int_st8_2[1] = dm_int_st7_2[2];
	// Bit 3
	full_adder FA840(.a(dm_int_st7_3[0]), .b(dm_int_st7_3[1]), .cin(dm_int_st7_3[2]), .s(dm_int_st8_3[1]), .cout(dm_int_st8_4[0]));
	// Bit 4
	full_adder FA841(.a(dm_int_st7_4[0]), .b(dm_int_st7_4[1]), .cin(dm_int_st7_4[2]), .s(dm_int_st8_4[1]), .cout(dm_int_st8_5[0]));
	// Bit 5
	full_adder FA842(.a(dm_int_st7_5[0]), .b(dm_int_st7_5[1]), .cin(dm_int_st7_5[2]), .s(dm_int_st8_5[1]), .cout(dm_int_st8_6[0]));
	// Bit 6
	full_adder FA843(.a(dm_int_st7_6[0]), .b(dm_int_st7_6[1]), .cin(dm_int_st7_6[2]), .s(dm_int_st8_6[1]), .cout(dm_int_st8_7[0]));
	// Bit 7
	full_adder FA844(.a(dm_int_st7_7[0]), .b(dm_int_st7_7[1]), .cin(dm_int_st7_7[2]), .s(dm_int_st8_7[1]), .cout(dm_int_st8_8[0]));
	// Bit 8
	full_adder FA845(.a(dm_int_st7_8[0]), .b(dm_int_st7_8[1]), .cin(dm_int_st7_8[2]), .s(dm_int_st8_8[1]), .cout(dm_int_st8_9[0]));
	// Bit 9
	full_adder FA846(.a(dm_int_st7_9[0]), .b(dm_int_st7_9[1]), .cin(dm_int_st7_9[2]), .s(dm_int_st8_9[1]), .cout(dm_int_st8_10[0]));
	// Bit 10
	full_adder FA847(.a(dm_int_st7_10[0]), .b(dm_int_st7_10[1]), .cin(dm_int_st7_10[2]), .s(dm_int_st8_10[1]), .cout(dm_int_st8_11[0]));
	// Bit 11
	full_adder FA848(.a(dm_int_st7_11[0]), .b(dm_int_st7_11[1]), .cin(dm_int_st7_11[2]), .s(dm_int_st8_11[1]), .cout(dm_int_st8_12[0]));
	// Bit 12
	full_adder FA849(.a(dm_int_st7_12[0]), .b(dm_int_st7_12[1]), .cin(dm_int_st7_12[2]), .s(dm_int_st8_12[1]), .cout(dm_int_st8_13[0]));
	// Bit 13
	full_adder FA850(.a(dm_int_st7_13[0]), .b(dm_int_st7_13[1]), .cin(dm_int_st7_13[2]), .s(dm_int_st8_13[1]), .cout(dm_int_st8_14[0]));
	// Bit 14
	full_adder FA851(.a(dm_int_st7_14[0]), .b(dm_int_st7_14[1]), .cin(dm_int_st7_14[2]), .s(dm_int_st8_14[1]), .cout(dm_int_st8_15[0]));
	// Bit 15
	full_adder FA852(.a(dm_int_st7_15[0]), .b(dm_int_st7_15[1]), .cin(dm_int_st7_15[2]), .s(dm_int_st8_15[1]), .cout(dm_int_st8_16[0]));
	// Bit 16
	full_adder FA853(.a(dm_int_st7_16[0]), .b(dm_int_st7_16[1]), .cin(dm_int_st7_16[2]), .s(dm_int_st8_16[1]), .cout(dm_int_st8_17[0]));
	// Bit 17
	full_adder FA854(.a(dm_int_st7_17[0]), .b(dm_int_st7_17[1]), .cin(dm_int_st7_17[2]), .s(dm_int_st8_17[1]), .cout(dm_int_st8_18[0]));
	// Bit 18
	full_adder FA855(.a(dm_int_st7_18[0]), .b(dm_int_st7_18[1]), .cin(dm_int_st7_18[2]), .s(dm_int_st8_18[1]), .cout(dm_int_st8_19[0]));
	// Bit 19
	full_adder FA856(.a(dm_int_st7_19[0]), .b(dm_int_st7_19[1]), .cin(dm_int_st7_19[2]), .s(dm_int_st8_19[1]), .cout(dm_int_st8_20[0]));
	// Bit 20
	full_adder FA857(.a(dm_int_st7_20[0]), .b(dm_int_st7_20[1]), .cin(dm_int_st7_20[2]), .s(dm_int_st8_20[1]), .cout(dm_int_st8_21[0]));
	// Bit 21
	full_adder FA858(.a(dm_int_st7_21[0]), .b(dm_int_st7_21[1]), .cin(dm_int_st7_21[2]), .s(dm_int_st8_21[1]), .cout(dm_int_st8_22[0]));
	// Bit 22
	full_adder FA859(.a(dm_int_st7_22[0]), .b(dm_int_st7_22[1]), .cin(dm_int_st7_22[2]), .s(dm_int_st8_22[1]), .cout(dm_int_st8_23[0]));
	// Bit 23
	full_adder FA860(.a(dm_int_st7_23[0]), .b(dm_int_st7_23[1]), .cin(dm_int_st7_23[2]), .s(dm_int_st8_23[1]), .cout(dm_int_st8_24[0]));
	// Bit 24
	full_adder FA861(.a(dm_int_st7_24[0]), .b(dm_int_st7_24[1]), .cin(dm_int_st7_24[2]), .s(dm_int_st8_24[1]), .cout(dm_int_st8_25[0]));
	// Bit 25
	full_adder FA862(.a(dm_int_st7_25[0]), .b(dm_int_st7_25[1]), .cin(dm_int_st7_25[2]), .s(dm_int_st8_25[1]), .cout(dm_int_st8_26[0]));
	// Bit 26
	full_adder FA863(.a(dm_int_st7_26[0]), .b(dm_int_st7_26[1]), .cin(dm_int_st7_26[2]), .s(dm_int_st8_26[1]), .cout(dm_int_st8_27[0]));
	// Bit 27
	full_adder FA864(.a(dm_int_st7_27[0]), .b(dm_int_st7_27[1]), .cin(dm_int_st7_27[2]), .s(dm_int_st8_27[1]), .cout(dm_int_st8_28[0]));
	// Bit 28
	full_adder FA865(.a(dm_int_st7_28[0]), .b(dm_int_st7_28[1]), .cin(dm_int_st7_28[2]), .s(dm_int_st8_28[1]), .cout(dm_int_st8_29[0]));
	// Bit 29
	full_adder FA866(.a(dm_int_st7_29[0]), .b(dm_int_st7_29[1]), .cin(dm_int_st7_29[2]), .s(dm_int_st8_29[1]), .cout(dm_int_st8_30[0]));
	// Bit 30
	full_adder FA867(.a(dm_int_st7_30[0]), .b(dm_int_st7_30[1]), .cin(dm_int_st7_30[2]), .s(dm_int_st8_30[1]), .cout(dm_int_st8_31[0]));
	// Bit 31
	full_adder FA868(.a(dm_int_st7_31[0]), .b(dm_int_st7_31[1]), .cin(dm_int_st7_31[2]), .s(dm_int_st8_31[1]), .cout(dm_int_st8_32[0]));
	// Bit 32
	full_adder FA869(.a(dm_int_st7_32[0]), .b(dm_int_st7_32[1]), .cin(dm_int_st7_32[2]), .s(dm_int_st8_32[1]), .cout(dm_int_st8_33[0]));
	// Bit 33
	full_adder FA870(.a(dm_int_st7_33[0]), .b(dm_int_st7_33[1]), .cin(dm_int_st7_33[2]), .s(dm_int_st8_33[1]), .cout(dm_int_st8_34[0]));
	// Bit 34
	full_adder FA871(.a(dm_int_st7_34[0]), .b(dm_int_st7_34[1]), .cin(dm_int_st7_34[2]), .s(dm_int_st8_34[1]), .cout(dm_int_st8_35[0]));
	// Bit 35
	full_adder FA872(.a(dm_int_st7_35[0]), .b(dm_int_st7_35[1]), .cin(dm_int_st7_35[2]), .s(dm_int_st8_35[1]), .cout(dm_int_st8_36[0]));
	// Bit 36
	full_adder FA873(.a(dm_int_st7_36[0]), .b(dm_int_st7_36[1]), .cin(dm_int_st7_36[2]), .s(dm_int_st8_36[1]), .cout(dm_int_st8_37[0]));
	// Bit 37
	full_adder FA874(.a(dm_int_st7_37[0]), .b(dm_int_st7_37[1]), .cin(dm_int_st7_37[2]), .s(dm_int_st8_37[1]), .cout(dm_int_st8_38[0]));
	// Bit 38
	full_adder FA875(.a(dm_int_st7_38[0]), .b(dm_int_st7_38[1]), .cin(dm_int_st7_38[2]), .s(dm_int_st8_38[1]), .cout(dm_int_st8_39[0]));
	// Bit 39
	full_adder FA876(.a(dm_int_st7_39[0]), .b(dm_int_st7_39[1]), .cin(dm_int_st7_39[2]), .s(dm_int_st8_39[1]), .cout(dm_int_st8_40[0]));
	// Bit 40
	full_adder FA877(.a(dm_int_st7_40[0]), .b(dm_int_st7_40[1]), .cin(dm_int_st7_40[2]), .s(dm_int_st8_40[1]), .cout(dm_int_st8_41[0]));
	// Bit 41
	full_adder FA878(.a(dm_int_st7_41[0]), .b(dm_int_st7_41[1]), .cin(dm_int_st7_41[2]), .s(dm_int_st8_41[1]), .cout(dm_int_st8_42[0]));
	// Bit 42
	full_adder FA879(.a(dm_int_st7_42[0]), .b(dm_int_st7_42[1]), .cin(dm_int_st7_42[2]), .s(dm_int_st8_42[1]), .cout(dm_int_st8_43[0]));
	// Bit 43
	full_adder FA880(.a(dm_int_st7_43[0]), .b(dm_int_st7_43[1]), .cin(dm_int_st7_43[2]), .s(dm_int_st8_43[1]), .cout(dm_int_st8_44[0]));
	// Bit 44
	full_adder FA881(.a(dm_int_st7_44[0]), .b(dm_int_st7_44[1]), .cin(dm_int_st7_44[2]), .s(dm_int_st8_44[1]), .cout(dm_int_st8_45[0]));
	// Bit 45
	full_adder FA882(.a(dm_int_st7_45[0]), .b(dm_int_st7_45[1]), .cin(dm_int_st7_45[2]), .s(dm_int_st8_45[1]), .cout(dm_int_st8_46[0]));
	// Bit 46
	full_adder FA883(.a(dm_int_st7_46[0]), .b(dm_int_st7_46[1]), .cin(dm_int_st7_46[2]), .s(dm_int_st8_46[1]), .cout(dm_int_st8_47[0]));
	// Bit 47
	full_adder FA884(.a(dm_int_st7_47[0]), .b(dm_int_st7_47[1]), .cin(dm_int_st7_47[2]), .s(dm_int_st8_47[1]), .cout(dm_int_st8_48[0]));
	// Bit 48
	full_adder FA885(.a(dm_int_st7_48[0]), .b(dm_int_st7_48[1]), .cin(dm_int_st7_48[2]), .s(dm_int_st8_48[1]), .cout(dm_int_st8_49[0]));
	// Bit 49
	full_adder FA886(.a(dm_int_st7_49[0]), .b(dm_int_st7_49[1]), .cin(dm_int_st7_49[2]), .s(dm_int_st8_49[1]), .cout(dm_int_st8_50[0]));
	// Bit 50
	full_adder FA887(.a(dm_int_st7_50[0]), .b(dm_int_st7_50[1]), .cin(dm_int_st7_50[2]), .s(dm_int_st8_50[1]), .cout(dm_int_st8_51[0]));
	// Bit 51
	full_adder FA888(.a(dm_int_st7_51[0]), .b(dm_int_st7_51[1]), .cin(dm_int_st7_51[2]), .s(dm_int_st8_51[1]), .cout(dm_int_st8_52[0]));
	// Bit 52
	full_adder FA889(.a(dm_int_st7_52[0]), .b(dm_int_st7_52[1]), .cin(dm_int_st7_52[2]), .s(dm_int_st8_52[1]), .cout(dm_int_st8_53[0]));
	// Bit 53
	full_adder FA890(.a(dm_int_st7_53[0]), .b(dm_int_st7_53[1]), .cin(dm_int_st7_53[2]), .s(dm_int_st8_53[1]), .cout(dm_int_st8_54[0]));
	// Bit 54
	full_adder FA891(.a(dm_int_st7_54[0]), .b(dm_int_st7_54[1]), .cin(dm_int_st7_54[2]), .s(dm_int_st8_54[1]), .cout(dm_int_st8_55[0]));
	// Bit 55
	full_adder FA892(.a(dm_int_st7_55[0]), .b(dm_int_st7_55[1]), .cin(dm_int_st7_55[2]), .s(dm_int_st8_55[1]), .cout(dm_int_st8_56[0]));
	// Bit 56
	full_adder FA893(.a(dm_int_st7_56[0]), .b(dm_int_st7_56[1]), .cin(dm_int_st7_56[2]), .s(dm_int_st8_56[1]), .cout(dm_int_st8_57[0]));
	// Bit 57
	full_adder FA894(.a(dm_int_st7_57[0]), .b(dm_int_st7_57[1]), .cin(dm_int_st7_57[2]), .s(dm_int_st8_57[1]), .cout(dm_int_st8_58[0]));
	// Bit 58
	full_adder FA895(.a(dm_int_st7_58[0]), .b(dm_int_st7_58[1]), .cin(dm_int_st7_58[2]), .s(dm_int_st8_58[1]), .cout(dm_int_st8_59[0]));
	// Bit 59
	full_adder FA896(.a(dm_int_st7_59[0]), .b(dm_int_st7_59[1]), .cin(dm_int_st7_59[2]), .s(dm_int_st8_59[1]), .cout(dm_int_st8_60[0]));
	// Bit 60
	full_adder FA897(.a(dm_int_st7_60[0]), .b(dm_int_st7_60[1]), .cin(dm_int_st7_60[2]), .s(dm_int_st8_60[1]), .cout(dm_int_st8_61[0]));
	// Bit 61
	full_adder FA898(.a(dm_int_st7_61[0]), .b(dm_int_st7_61[1]), .cin(dm_int_st7_61[2]), .s(dm_int_st8_61[1]), .cout(dm_int_st8_62[0]));
	// Bit 62
	assign dm_int_st8_62[1] = dm_int_st7_62[0];

	// Adder Stage
	wire [63:0] cla_in_a, cla_in_b, sum;
	wire ovf;
	assign cla_in_a[0] = dm_int_st8_0[0];
	assign cla_in_b[0] = 1'b0;
	assign cla_in_a[1] = dm_int_st8_1[0];
	assign cla_in_b[1] = dm_int_st8_1[1];
	assign cla_in_a[2] = dm_int_st8_2[0];
	assign cla_in_b[2] = dm_int_st8_2[1];
	assign cla_in_a[3] = dm_int_st8_3[0];
	assign cla_in_b[3] = dm_int_st8_3[1];
	assign cla_in_a[4] = dm_int_st8_4[0];
	assign cla_in_b[4] = dm_int_st8_4[1];
	assign cla_in_a[5] = dm_int_st8_5[0];
	assign cla_in_b[5] = dm_int_st8_5[1];
	assign cla_in_a[6] = dm_int_st8_6[0];
	assign cla_in_b[6] = dm_int_st8_6[1];
	assign cla_in_a[7] = dm_int_st8_7[0];
	assign cla_in_b[7] = dm_int_st8_7[1];
	assign cla_in_a[8] = dm_int_st8_8[0];
	assign cla_in_b[8] = dm_int_st8_8[1];
	assign cla_in_a[9] = dm_int_st8_9[0];
	assign cla_in_b[9] = dm_int_st8_9[1];
	assign cla_in_a[10] = dm_int_st8_10[0];
	assign cla_in_b[10] = dm_int_st8_10[1];
	assign cla_in_a[11] = dm_int_st8_11[0];
	assign cla_in_b[11] = dm_int_st8_11[1];
	assign cla_in_a[12] = dm_int_st8_12[0];
	assign cla_in_b[12] = dm_int_st8_12[1];
	assign cla_in_a[13] = dm_int_st8_13[0];
	assign cla_in_b[13] = dm_int_st8_13[1];
	assign cla_in_a[14] = dm_int_st8_14[0];
	assign cla_in_b[14] = dm_int_st8_14[1];
	assign cla_in_a[15] = dm_int_st8_15[0];
	assign cla_in_b[15] = dm_int_st8_15[1];
	assign cla_in_a[16] = dm_int_st8_16[0];
	assign cla_in_b[16] = dm_int_st8_16[1];
	assign cla_in_a[17] = dm_int_st8_17[0];
	assign cla_in_b[17] = dm_int_st8_17[1];
	assign cla_in_a[18] = dm_int_st8_18[0];
	assign cla_in_b[18] = dm_int_st8_18[1];
	assign cla_in_a[19] = dm_int_st8_19[0];
	assign cla_in_b[19] = dm_int_st8_19[1];
	assign cla_in_a[20] = dm_int_st8_20[0];
	assign cla_in_b[20] = dm_int_st8_20[1];
	assign cla_in_a[21] = dm_int_st8_21[0];
	assign cla_in_b[21] = dm_int_st8_21[1];
	assign cla_in_a[22] = dm_int_st8_22[0];
	assign cla_in_b[22] = dm_int_st8_22[1];
	assign cla_in_a[23] = dm_int_st8_23[0];
	assign cla_in_b[23] = dm_int_st8_23[1];
	assign cla_in_a[24] = dm_int_st8_24[0];
	assign cla_in_b[24] = dm_int_st8_24[1];
	assign cla_in_a[25] = dm_int_st8_25[0];
	assign cla_in_b[25] = dm_int_st8_25[1];
	assign cla_in_a[26] = dm_int_st8_26[0];
	assign cla_in_b[26] = dm_int_st8_26[1];
	assign cla_in_a[27] = dm_int_st8_27[0];
	assign cla_in_b[27] = dm_int_st8_27[1];
	assign cla_in_a[28] = dm_int_st8_28[0];
	assign cla_in_b[28] = dm_int_st8_28[1];
	assign cla_in_a[29] = dm_int_st8_29[0];
	assign cla_in_b[29] = dm_int_st8_29[1];
	assign cla_in_a[30] = dm_int_st8_30[0];
	assign cla_in_b[30] = dm_int_st8_30[1];
	assign cla_in_a[31] = dm_int_st8_31[0];
	assign cla_in_b[31] = dm_int_st8_31[1];
	assign cla_in_a[32] = dm_int_st8_32[0];
	assign cla_in_b[32] = dm_int_st8_32[1];
	assign cla_in_a[33] = dm_int_st8_33[0];
	assign cla_in_b[33] = dm_int_st8_33[1];
	assign cla_in_a[34] = dm_int_st8_34[0];
	assign cla_in_b[34] = dm_int_st8_34[1];
	assign cla_in_a[35] = dm_int_st8_35[0];
	assign cla_in_b[35] = dm_int_st8_35[1];
	assign cla_in_a[36] = dm_int_st8_36[0];
	assign cla_in_b[36] = dm_int_st8_36[1];
	assign cla_in_a[37] = dm_int_st8_37[0];
	assign cla_in_b[37] = dm_int_st8_37[1];
	assign cla_in_a[38] = dm_int_st8_38[0];
	assign cla_in_b[38] = dm_int_st8_38[1];
	assign cla_in_a[39] = dm_int_st8_39[0];
	assign cla_in_b[39] = dm_int_st8_39[1];
	assign cla_in_a[40] = dm_int_st8_40[0];
	assign cla_in_b[40] = dm_int_st8_40[1];
	assign cla_in_a[41] = dm_int_st8_41[0];
	assign cla_in_b[41] = dm_int_st8_41[1];
	assign cla_in_a[42] = dm_int_st8_42[0];
	assign cla_in_b[42] = dm_int_st8_42[1];
	assign cla_in_a[43] = dm_int_st8_43[0];
	assign cla_in_b[43] = dm_int_st8_43[1];
	assign cla_in_a[44] = dm_int_st8_44[0];
	assign cla_in_b[44] = dm_int_st8_44[1];
	assign cla_in_a[45] = dm_int_st8_45[0];
	assign cla_in_b[45] = dm_int_st8_45[1];
	assign cla_in_a[46] = dm_int_st8_46[0];
	assign cla_in_b[46] = dm_int_st8_46[1];
	assign cla_in_a[47] = dm_int_st8_47[0];
	assign cla_in_b[47] = dm_int_st8_47[1];
	assign cla_in_a[48] = dm_int_st8_48[0];
	assign cla_in_b[48] = dm_int_st8_48[1];
	assign cla_in_a[49] = dm_int_st8_49[0];
	assign cla_in_b[49] = dm_int_st8_49[1];
	assign cla_in_a[50] = dm_int_st8_50[0];
	assign cla_in_b[50] = dm_int_st8_50[1];
	assign cla_in_a[51] = dm_int_st8_51[0];
	assign cla_in_b[51] = dm_int_st8_51[1];
	assign cla_in_a[52] = dm_int_st8_52[0];
	assign cla_in_b[52] = dm_int_st8_52[1];
	assign cla_in_a[53] = dm_int_st8_53[0];
	assign cla_in_b[53] = dm_int_st8_53[1];
	assign cla_in_a[54] = dm_int_st8_54[0];
	assign cla_in_b[54] = dm_int_st8_54[1];
	assign cla_in_a[55] = dm_int_st8_55[0];
	assign cla_in_b[55] = dm_int_st8_55[1];
	assign cla_in_a[56] = dm_int_st8_56[0];
	assign cla_in_b[56] = dm_int_st8_56[1];
	assign cla_in_a[57] = dm_int_st8_57[0];
	assign cla_in_b[57] = dm_int_st8_57[1];
	assign cla_in_a[58] = dm_int_st8_58[0];
	assign cla_in_b[58] = dm_int_st8_58[1];
	assign cla_in_a[59] = dm_int_st8_59[0];
	assign cla_in_b[59] = dm_int_st8_59[1];
	assign cla_in_a[60] = dm_int_st8_60[0];
	assign cla_in_b[60] = dm_int_st8_60[1];
	assign cla_in_a[61] = dm_int_st8_61[0];
	assign cla_in_b[61] = dm_int_st8_61[1];
	assign cla_in_a[62] = dm_int_st8_62[0];
	assign cla_in_b[62] = dm_int_st8_62[1];
	assign cla_in_a[63] = 1'b0;
	assign cla_in_b[63] = 1'b0;
	cla_64bit CLA(clk, cla_in_a, cla_in_b, 1'b0, sum, ovf);

	assign out_overflow = sum[61];
	assign out_s[`FXP32S_MAG] = sum[60:30] | {`FXP32S_WIDTH-1{out_overflow}};
	assign out_s[`FXP32S_SIGN] = neg_out;

endmodule
